--! Standard libraries
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--! User packages
use work.tf_pkg.all;
use work.memUtil_pkg.all;

entity SectorProcessor is
  port(
    clk        : in std_logic;
    reset      : in std_logic;
    IR_start  : in std_logic;
    IR_bx_in : in std_logic_vector(2 downto 0);
    TP_bx_out_merged : out std_logic_vector(2 downto 0);
    TP_bx_out : out std_logic_vector(2 downto 0);
    TP_bx_out_vld : out std_logic;
    TP_done   : out std_logic;
    DL_PS10G_1_A_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_1_A_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_1_A_link_read          : out t_DL_39_1b;
    DL_PS10G_1_B_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_1_B_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_1_B_link_read          : out t_DL_39_1b;
    DL_PS10G_2_A_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_2_A_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_2_A_link_read          : out t_DL_39_1b;
    DL_PS10G_2_B_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_2_B_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_2_B_link_read          : out t_DL_39_1b;
    DL_PS10G_3_A_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_3_A_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_3_A_link_read          : out t_DL_39_1b;
    DL_PS10G_3_B_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_3_B_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_3_B_link_read          : out t_DL_39_1b;
    DL_PS10G_4_A_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_4_A_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_4_A_link_read          : out t_DL_39_1b;
    DL_PS10G_4_B_link_AV_dout       : in t_DL_39_DATA;
    DL_PS10G_4_B_link_empty_neg     : in t_DL_39_1b;
    DL_PS10G_4_B_link_read          : out t_DL_39_1b;
    DL_PS_1_A_link_AV_dout       : in t_DL_39_DATA;
    DL_PS_1_A_link_empty_neg     : in t_DL_39_1b;
    DL_PS_1_A_link_read          : out t_DL_39_1b;
    DL_PS_1_B_link_AV_dout       : in t_DL_39_DATA;
    DL_PS_1_B_link_empty_neg     : in t_DL_39_1b;
    DL_PS_1_B_link_read          : out t_DL_39_1b;
    DL_PS_2_A_link_AV_dout       : in t_DL_39_DATA;
    DL_PS_2_A_link_empty_neg     : in t_DL_39_1b;
    DL_PS_2_A_link_read          : out t_DL_39_1b;
    DL_PS_2_B_link_AV_dout       : in t_DL_39_DATA;
    DL_PS_2_B_link_empty_neg     : in t_DL_39_1b;
    DL_PS_2_B_link_read          : out t_DL_39_1b;
    DL_negPS10G_1_A_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_1_A_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_1_A_link_read          : out t_DL_39_1b;
    DL_negPS10G_1_B_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_1_B_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_1_B_link_read          : out t_DL_39_1b;
    DL_negPS10G_2_A_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_2_A_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_2_A_link_read          : out t_DL_39_1b;
    DL_negPS10G_2_B_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_2_B_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_2_B_link_read          : out t_DL_39_1b;
    DL_negPS10G_3_A_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_3_A_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_3_A_link_read          : out t_DL_39_1b;
    DL_negPS10G_3_B_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_3_B_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_3_B_link_read          : out t_DL_39_1b;
    DL_negPS10G_4_A_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_4_A_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_4_A_link_read          : out t_DL_39_1b;
    DL_negPS10G_4_B_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS10G_4_B_link_empty_neg     : in t_DL_39_1b;
    DL_negPS10G_4_B_link_read          : out t_DL_39_1b;
    DL_negPS_1_A_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS_1_A_link_empty_neg     : in t_DL_39_1b;
    DL_negPS_1_A_link_read          : out t_DL_39_1b;
    DL_negPS_1_B_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS_1_B_link_empty_neg     : in t_DL_39_1b;
    DL_negPS_1_B_link_read          : out t_DL_39_1b;
    DL_negPS_2_A_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS_2_A_link_empty_neg     : in t_DL_39_1b;
    DL_negPS_2_A_link_read          : out t_DL_39_1b;
    DL_negPS_2_B_link_AV_dout       : in t_DL_39_DATA;
    DL_negPS_2_B_link_empty_neg     : in t_DL_39_1b;
    DL_negPS_2_B_link_read          : out t_DL_39_1b;
    DL_twoS_1_A_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_1_A_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_1_A_link_read          : out t_DL_39_1b;
    DL_twoS_1_B_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_1_B_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_1_B_link_read          : out t_DL_39_1b;
    DL_twoS_2_A_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_2_A_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_2_A_link_read          : out t_DL_39_1b;
    DL_twoS_2_B_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_2_B_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_2_B_link_read          : out t_DL_39_1b;
    DL_twoS_3_A_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_3_A_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_3_A_link_read          : out t_DL_39_1b;
    DL_twoS_3_B_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_3_B_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_3_B_link_read          : out t_DL_39_1b;
    DL_twoS_4_A_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_4_A_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_4_A_link_read          : out t_DL_39_1b;
    DL_twoS_4_B_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_4_B_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_4_B_link_read          : out t_DL_39_1b;
    DL_twoS_5_A_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_5_A_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_5_A_link_read          : out t_DL_39_1b;
    DL_twoS_5_B_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_5_B_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_5_B_link_read          : out t_DL_39_1b;
    DL_twoS_6_A_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_6_A_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_6_A_link_read          : out t_DL_39_1b;
    DL_twoS_6_B_link_AV_dout       : in t_DL_39_DATA;
    DL_twoS_6_B_link_empty_neg     : in t_DL_39_1b;
    DL_twoS_6_B_link_read          : out t_DL_39_1b;
    DL_neg2S_1_A_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_1_A_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_1_A_link_read          : out t_DL_39_1b;
    DL_neg2S_1_B_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_1_B_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_1_B_link_read          : out t_DL_39_1b;
    DL_neg2S_2_A_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_2_A_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_2_A_link_read          : out t_DL_39_1b;
    DL_neg2S_2_B_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_2_B_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_2_B_link_read          : out t_DL_39_1b;
    DL_neg2S_3_A_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_3_A_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_3_A_link_read          : out t_DL_39_1b;
    DL_neg2S_3_B_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_3_B_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_3_B_link_read          : out t_DL_39_1b;
    DL_neg2S_4_A_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_4_A_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_4_A_link_read          : out t_DL_39_1b;
    DL_neg2S_4_B_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_4_B_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_4_B_link_read          : out t_DL_39_1b;
    DL_neg2S_5_A_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_5_A_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_5_A_link_read          : out t_DL_39_1b;
    DL_neg2S_5_B_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_5_B_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_5_B_link_read          : out t_DL_39_1b;
    DL_neg2S_6_A_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_6_A_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_6_A_link_read          : out t_DL_39_1b;
    DL_neg2S_6_B_link_AV_dout       : in t_DL_39_DATA;
    DL_neg2S_6_B_link_empty_neg     : in t_DL_39_1b;
    DL_neg2S_6_B_link_read          : out t_DL_39_1b;
    --AS_L1PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L1PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L1PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L1PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L1PHIEn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L1PHIFn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L1PHIGn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L1PHIHn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L2PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L2PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L2PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L2PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L3PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L3PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L3PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L3PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L4PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L4PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L4PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L4PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L5PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L5PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L5PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L5PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L6PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L6PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L6PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_L6PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D1PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D1PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D1PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D1PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D2PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D2PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D2PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D2PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D3PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D3PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D3PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D3PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D4PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D4PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D4PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D4PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D5PHIAn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D5PHIBn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D5PHICn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --AS_D5PHIDn1_stream_V_dout : out std_logic_vector(36 downto 0);
    --MPAR_L1L2ABC_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L1L2DE_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L1L2F_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L1L2G_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L1L2HI_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L1L2JKL_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L2L3ABCD_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L3L4AB_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L3L4CD_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L5L6ABCD_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_D1D2ABCD_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_D3D4ABCD_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L1D1ABCD_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L1D1EFGH_stream_V_dout : out std_logic_vector(75 downto 0);
    --MPAR_L2D1ABCD_stream_V_dout : out std_logic_vector(75 downto 0)



    AS_D1PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_D1PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_D1PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_D1PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_D2PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_D2PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_D2PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_D2PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_D3PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_D3PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_D3PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_D3PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_D4PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_D4PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_D4PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_D4PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_D5PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_D5PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_D5PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_D5PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHIEn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHIFn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHIGn1_V_readaddr : in t_AS_36_ADDR;
    AS_L1PHIHn1_V_readaddr : in t_AS_36_ADDR;
    AS_L2PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_L2PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_L2PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_L2PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_L3PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_L3PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_L3PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_L3PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_L4PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_L4PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_L4PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_L4PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_L5PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_L5PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_L5PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_L5PHIDn1_V_readaddr : in t_AS_36_ADDR;
    AS_L6PHIAn1_V_readaddr : in t_AS_36_ADDR;
    AS_L6PHIBn1_V_readaddr : in t_AS_36_ADDR;
    AS_L6PHICn1_V_readaddr : in t_AS_36_ADDR;
    AS_L6PHIDn1_V_readaddr : in t_AS_36_ADDR;
    TPAR_D1D2A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_D1D2B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_D1D2C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_D1D2D_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_D3D4A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_D3D4B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_D3D4C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_D3D4D_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1D_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1E_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1F_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1G_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1D1H_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2D_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2E_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2F_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2G_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2H_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2I_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2J_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2K_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L1L2L_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2D1A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2D1B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2D1C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2D1D_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2L3A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2L3B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2L3C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L2L3D_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L3L4A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L3L4B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L3L4C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L3L4D_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L5L6A_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L5L6B_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L5L6C_V_readaddr : in t_TPAR_73_ADDR;
    TPAR_L5L6D_V_readaddr : in t_TPAR_73_ADDR;

    AS_D1PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D1PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_D1PHIAn1_bx_vld : out std_logic;
    AS_D1PHIAn1_V_dout : out t_AS_36_DATA;
    AS_D1PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D1PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_D1PHIBn1_bx_vld : out std_logic;
    AS_D1PHIBn1_V_dout : out t_AS_36_DATA;
    AS_D1PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D1PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_D1PHICn1_bx_vld : out std_logic;
    AS_D1PHICn1_V_dout : out t_AS_36_DATA;
    AS_D1PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D1PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_D1PHIDn1_bx_vld : out std_logic;
    AS_D1PHIDn1_V_dout : out t_AS_36_DATA;
    AS_D2PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D2PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_D2PHIAn1_bx_vld : out std_logic;
    AS_D2PHIAn1_V_dout : out t_AS_36_DATA;
    AS_D2PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D2PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_D2PHIBn1_bx_vld : out std_logic;
    AS_D2PHIBn1_V_dout : out t_AS_36_DATA;
    AS_D2PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D2PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_D2PHICn1_bx_vld : out std_logic;
    AS_D2PHICn1_V_dout : out t_AS_36_DATA;
    AS_D2PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D2PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_D2PHIDn1_bx_vld : out std_logic;
    AS_D2PHIDn1_V_dout : out t_AS_36_DATA;
    AS_D3PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D3PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_D3PHIAn1_bx_vld : out std_logic;
    AS_D3PHIAn1_V_dout : out t_AS_36_DATA;
    AS_D3PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D3PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_D3PHIBn1_bx_vld : out std_logic;
    AS_D3PHIBn1_V_dout : out t_AS_36_DATA;
    AS_D3PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D3PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_D3PHICn1_bx_vld : out std_logic;
    AS_D3PHICn1_V_dout : out t_AS_36_DATA;
    AS_D3PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D3PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_D3PHIDn1_bx_vld : out std_logic;
    AS_D3PHIDn1_V_dout : out t_AS_36_DATA;
    AS_D4PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D4PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_D4PHIAn1_bx_vld : out std_logic;
    AS_D4PHIAn1_V_dout : out t_AS_36_DATA;
    AS_D4PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D4PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_D4PHIBn1_bx_vld : out std_logic;
    AS_D4PHIBn1_V_dout : out t_AS_36_DATA;
    AS_D4PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D4PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_D4PHICn1_bx_vld : out std_logic;
    AS_D4PHICn1_V_dout : out t_AS_36_DATA;
    AS_D4PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D4PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_D4PHIDn1_bx_vld : out std_logic;
    AS_D4PHIDn1_V_dout : out t_AS_36_DATA;
    AS_D5PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D5PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_D5PHIAn1_bx_vld : out std_logic;
    AS_D5PHIAn1_V_dout : out t_AS_36_DATA;
    AS_D5PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D5PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_D5PHIBn1_bx_vld : out std_logic;
    AS_D5PHIBn1_V_dout : out t_AS_36_DATA;
    AS_D5PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D5PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_D5PHICn1_bx_vld : out std_logic;
    AS_D5PHICn1_V_dout : out t_AS_36_DATA;
    AS_D5PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_D5PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_D5PHIDn1_bx_vld : out std_logic;
    AS_D5PHIDn1_V_dout : out t_AS_36_DATA;
    AS_L1PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHIAn1_bx_vld : out std_logic;
    AS_L1PHIAn1_V_dout : out t_AS_36_DATA;
    AS_L1PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHIBn1_bx_vld : out std_logic;
    AS_L1PHIBn1_V_dout : out t_AS_36_DATA;
    AS_L1PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHICn1_bx_vld : out std_logic;
    AS_L1PHICn1_V_dout : out t_AS_36_DATA;
    AS_L1PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHIDn1_bx_vld : out std_logic;
    AS_L1PHIDn1_V_dout : out t_AS_36_DATA;
    AS_L1PHIEn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHIEn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHIEn1_bx_vld : out std_logic;
    AS_L1PHIEn1_V_dout : out t_AS_36_DATA;
    AS_L1PHIFn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHIFn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHIFn1_bx_vld : out std_logic;
    AS_L1PHIFn1_V_dout : out t_AS_36_DATA;
    AS_L1PHIGn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHIGn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHIGn1_bx_vld : out std_logic;
    AS_L1PHIGn1_V_dout : out t_AS_36_DATA;
    AS_L1PHIHn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L1PHIHn1_bx : out std_logic_vector(2 downto 0);
    AS_L1PHIHn1_bx_vld : out std_logic;
    AS_L1PHIHn1_V_dout : out t_AS_36_DATA;
    AS_L2PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L2PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_L2PHIAn1_bx_vld : out std_logic;
    AS_L2PHIAn1_V_dout : out t_AS_36_DATA;
    AS_L2PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L2PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_L2PHIBn1_bx_vld : out std_logic;
    AS_L2PHIBn1_V_dout : out t_AS_36_DATA;
    AS_L2PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L2PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_L2PHICn1_bx_vld : out std_logic;
    AS_L2PHICn1_V_dout : out t_AS_36_DATA;
    AS_L2PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L2PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_L2PHIDn1_bx_vld : out std_logic;
    AS_L2PHIDn1_V_dout : out t_AS_36_DATA;
    AS_L3PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L3PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_L3PHIAn1_bx_vld : out std_logic;
    AS_L3PHIAn1_V_dout : out t_AS_36_DATA;
    AS_L3PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L3PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_L3PHIBn1_bx_vld : out std_logic;
    AS_L3PHIBn1_V_dout : out t_AS_36_DATA;
    AS_L3PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L3PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_L3PHICn1_bx_vld : out std_logic;
    AS_L3PHICn1_V_dout : out t_AS_36_DATA;
    AS_L3PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L3PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_L3PHIDn1_bx_vld : out std_logic;
    AS_L3PHIDn1_V_dout : out t_AS_36_DATA;
    AS_L4PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L4PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_L4PHIAn1_bx_vld : out std_logic;
    AS_L4PHIAn1_V_dout : out t_AS_36_DATA;
    AS_L4PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L4PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_L4PHIBn1_bx_vld : out std_logic;
    AS_L4PHIBn1_V_dout : out t_AS_36_DATA;
    AS_L4PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L4PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_L4PHICn1_bx_vld : out std_logic;
    AS_L4PHICn1_V_dout : out t_AS_36_DATA;
    AS_L4PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L4PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_L4PHIDn1_bx_vld : out std_logic;
    AS_L4PHIDn1_V_dout : out t_AS_36_DATA;
    AS_L5PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L5PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_L5PHIAn1_bx_vld : out std_logic;
    AS_L5PHIAn1_V_dout : out t_AS_36_DATA;
    AS_L5PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L5PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_L5PHIBn1_bx_vld : out std_logic;
    AS_L5PHIBn1_V_dout : out t_AS_36_DATA;
    AS_L5PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L5PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_L5PHICn1_bx_vld : out std_logic;
    AS_L5PHICn1_V_dout : out t_AS_36_DATA;
    AS_L5PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L5PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_L5PHIDn1_bx_vld : out std_logic;
    AS_L5PHIDn1_V_dout : out t_AS_36_DATA;
    AS_L6PHIAn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L6PHIAn1_bx : out std_logic_vector(2 downto 0);
    AS_L6PHIAn1_bx_vld : out std_logic;
    AS_L6PHIAn1_V_dout : out t_AS_36_DATA;
    AS_L6PHIBn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L6PHIBn1_bx : out std_logic_vector(2 downto 0);
    AS_L6PHIBn1_bx_vld : out std_logic;
    AS_L6PHIBn1_V_dout : out t_AS_36_DATA;
    AS_L6PHICn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L6PHICn1_bx : out std_logic_vector(2 downto 0);
    AS_L6PHICn1_bx_vld : out std_logic;
    AS_L6PHICn1_V_dout : out t_AS_36_DATA;
    AS_L6PHIDn1_AV_dout_nent : out t_AS_36_NENT;
    AS_L6PHIDn1_bx : out std_logic_vector(2 downto 0);
    AS_L6PHIDn1_bx_vld : out std_logic;
    AS_L6PHIDn1_V_dout : out t_AS_36_DATA;
    TPAR_D1D2A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARD1D2ABCD_bx : out std_logic_vector(2 downto 0);
    TPARD1D2ABCD_bx_vld : out std_logic;
    TPAR_D1D2A_V_dout : out t_TPAR_73_DATA;
    TPAR_D1D2B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_D1D2B_V_dout : out t_TPAR_73_DATA;
    TPAR_D1D2C_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_D1D2C_V_dout : out t_TPAR_73_DATA;
    TPAR_D1D2D_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_D1D2D_V_dout : out t_TPAR_73_DATA;
    TPAR_D3D4A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARD3D4ABCD_bx : out std_logic_vector(2 downto 0);
    TPARD3D4ABCD_bx_vld : out std_logic;
    TPAR_D3D4A_V_dout : out t_TPAR_73_DATA;
    TPAR_D3D4B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_D3D4B_V_dout : out t_TPAR_73_DATA;
    TPAR_D3D4C_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_D3D4C_V_dout : out t_TPAR_73_DATA;
    TPAR_D3D4D_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_D3D4D_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1D1ABCD_bx : out std_logic_vector(2 downto 0);
    TPARL1D1ABCD_bx_vld : out std_logic;
    TPAR_L1D1A_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1D1B_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1C_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1D1C_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1D_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1D1D_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1E_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1D1EFGH_bx : out std_logic_vector(2 downto 0);
    TPARL1D1EFGH_bx_vld : out std_logic;
    TPAR_L1D1E_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1F_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1D1F_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1G_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1D1G_V_dout : out t_TPAR_73_DATA;
    TPAR_L1D1H_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1D1H_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1L2ABC_bx : out std_logic_vector(2 downto 0);
    TPARL1L2ABC_bx_vld : out std_logic;
    TPAR_L1L2A_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1L2B_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2C_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1L2C_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2D_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1L2DE_bx : out std_logic_vector(2 downto 0);
    TPARL1L2DE_bx_vld : out std_logic;
    TPAR_L1L2D_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2E_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1L2E_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2F_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1L2F_bx : out std_logic_vector(2 downto 0);
    TPARL1L2F_bx_vld : out std_logic;
    TPAR_L1L2F_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2G_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1L2G_bx : out std_logic_vector(2 downto 0);
    TPARL1L2G_bx_vld : out std_logic;
    TPAR_L1L2G_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2H_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1L2HI_bx : out std_logic_vector(2 downto 0);
    TPARL1L2HI_bx_vld : out std_logic;
    TPAR_L1L2H_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2I_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1L2I_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2J_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL1L2JKL_bx : out std_logic_vector(2 downto 0);
    TPARL1L2JKL_bx_vld : out std_logic;
    TPAR_L1L2J_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2K_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1L2K_V_dout : out t_TPAR_73_DATA;
    TPAR_L1L2L_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L1L2L_V_dout : out t_TPAR_73_DATA;
    TPAR_L2D1A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL2D1ABCD_bx : out std_logic_vector(2 downto 0);
    TPARL2D1ABCD_bx_vld : out std_logic;
    TPAR_L2D1A_V_dout : out t_TPAR_73_DATA;
    TPAR_L2D1B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L2D1B_V_dout : out t_TPAR_73_DATA;
    TPAR_L2D1C_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L2D1C_V_dout : out t_TPAR_73_DATA;
    TPAR_L2D1D_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L2D1D_V_dout : out t_TPAR_73_DATA;
    TPAR_L2L3A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL2L3ABCD_bx : out std_logic_vector(2 downto 0);
    TPARL2L3ABCD_bx_vld : out std_logic;
    TPAR_L2L3A_V_dout : out t_TPAR_73_DATA;
    TPAR_L2L3B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L2L3B_V_dout : out t_TPAR_73_DATA;
    TPAR_L2L3C_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L2L3C_V_dout : out t_TPAR_73_DATA;
    TPAR_L2L3D_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L2L3D_V_dout : out t_TPAR_73_DATA;
    TPAR_L3L4A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL3L4AB_bx : out std_logic_vector(2 downto 0);
    TPARL3L4AB_bx_vld : out std_logic;
    TPAR_L3L4A_V_dout : out t_TPAR_73_DATA;
    TPAR_L3L4B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L3L4B_V_dout : out t_TPAR_73_DATA;
    TPAR_L3L4C_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL3L4CD_bx : out std_logic_vector(2 downto 0);
    TPARL3L4CD_bx_vld : out std_logic;
    TPAR_L3L4C_V_dout : out t_TPAR_73_DATA;
    TPAR_L3L4D_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L3L4D_V_dout : out t_TPAR_73_DATA;
    TPAR_L5L6A_AV_dout_nent : out t_TPAR_73_NENT;
    TPARL5L6ABCD_bx : out std_logic_vector(2 downto 0);
    TPARL5L6ABCD_bx_vld : out std_logic;
    TPAR_L5L6A_V_dout : out t_TPAR_73_DATA;
    TPAR_L5L6B_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L5L6B_V_dout : out t_TPAR_73_DATA;
    TPAR_L5L6C_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L5L6C_V_dout : out t_TPAR_73_DATA;
    TPAR_L5L6D_AV_dout_nent : out t_TPAR_73_NENT;
    TPAR_L5L6D_V_dout : out t_TPAR_73_DATA
  );
end SectorProcessor;

architecture rtl of SectorProcessor is

  signal IL_L1PHIA_PS10G_1_A_start                   : std_logic;
  signal IL_L1PHIA_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIA_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIA_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIA_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_L1PHIA_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIA_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_L1PHIA_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIA_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIA_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIA_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIB_PS10G_1_A_start                   : std_logic;
  signal IL_L1PHIB_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIB_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIB_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIB_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_L1PHIB_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIB_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_L1PHIB_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIB_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIB_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIB_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIC_PS10G_1_A_start                   : std_logic;
  signal IL_L1PHIC_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIC_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIC_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIC_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_L1PHIC_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIC_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_L1PHIC_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIC_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIC_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIC_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHID_PS10G_1_A_start                   : std_logic;
  signal IL_L1PHID_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHID_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_L1PHID_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHID_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIE_PS10G_1_A_start                   : std_logic;
  signal IL_L1PHIE_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIE_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_L1PHIE_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIE_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIG_PS10G_1_B_start                   : std_logic;
  signal IL_L1PHIG_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIG_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIG_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIG_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_L1PHIG_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIG_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_L1PHIG_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIG_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIG_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIG_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIH_PS10G_1_B_start                   : std_logic;
  signal IL_L1PHIH_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIH_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIH_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIH_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_L1PHIH_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIH_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_L1PHIH_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIH_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIH_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIH_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIA_PS10G_1_A_start                   : std_logic;
  signal IL_D1PHIA_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIA_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIA_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIA_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D1PHIA_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIA_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D1PHIA_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIA_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIA_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIA_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_PS10G_1_A_start                   : std_logic;
  signal IL_D1PHIB_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_PS10G_1_B_start                   : std_logic;
  signal IL_D1PHIB_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_PS10G_1_A_start                   : std_logic;
  signal IL_D1PHIC_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_PS10G_1_B_start                   : std_logic;
  signal IL_D1PHIC_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHID_PS10G_1_B_start                   : std_logic;
  signal IL_D1PHID_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHID_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHID_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHID_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D1PHID_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHID_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D1PHID_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHID_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHID_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHID_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIA_PS10G_1_A_start                   : std_logic;
  signal IL_D3PHIA_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIA_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIA_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIA_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D3PHIA_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIA_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D3PHIA_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIA_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIA_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIA_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_PS10G_1_A_start                   : std_logic;
  signal IL_D3PHIB_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_PS10G_1_B_start                   : std_logic;
  signal IL_D3PHIB_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_PS10G_1_A_start                   : std_logic;
  signal IL_D3PHIC_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_PS10G_1_B_start                   : std_logic;
  signal IL_D3PHIC_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHID_PS10G_1_B_start                   : std_logic;
  signal IL_D3PHID_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHID_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHID_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHID_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D3PHID_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHID_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D3PHID_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHID_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHID_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHID_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIA_PS10G_1_A_start                   : std_logic;
  signal IL_D5PHIA_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIA_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIA_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIA_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D5PHIA_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIA_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D5PHIA_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIA_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIA_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIA_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_PS10G_1_A_start                   : std_logic;
  signal IL_D5PHIB_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_PS10G_1_B_start                   : std_logic;
  signal IL_D5PHIB_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_PS10G_1_A_start                   : std_logic;
  signal IL_D5PHIC_PS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_PS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_PS10G_1_B_start                   : std_logic;
  signal IL_D5PHIC_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHID_PS10G_1_B_start                   : std_logic;
  signal IL_D5PHID_PS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHID_PS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHID_PS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHID_PS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D5PHID_PS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHID_PS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D5PHID_PS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHID_PS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHID_PS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHID_PS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIA_PS10G_2_A_start                   : std_logic;
  signal IL_L1PHIA_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIA_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIA_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIA_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIA_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIA_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIA_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIA_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIA_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIA_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIB_PS10G_2_A_start                   : std_logic;
  signal IL_L1PHIB_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIB_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIB_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIB_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIB_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIB_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIB_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIB_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIB_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIB_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIC_PS10G_2_A_start                   : std_logic;
  signal IL_L1PHIC_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIC_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIC_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIC_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIC_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIC_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIC_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIC_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIC_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIC_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHID_PS10G_2_A_start                   : std_logic;
  signal IL_L1PHID_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHID_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHID_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHID_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHID_PS10G_2_B_start                   : std_logic;
  signal IL_L1PHID_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHID_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHID_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHID_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHID_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHID_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIE_PS10G_2_A_start                   : std_logic;
  signal IL_L1PHIE_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIE_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIE_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIE_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIE_PS10G_2_B_start                   : std_logic;
  signal IL_L1PHIE_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIE_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIE_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIE_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIE_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIE_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIF_PS10G_2_B_start                   : std_logic;
  signal IL_L1PHIF_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIF_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIF_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIF_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIF_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIF_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIF_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIF_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIF_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIF_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIG_PS10G_2_B_start                   : std_logic;
  signal IL_L1PHIG_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIG_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIG_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIG_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIG_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIG_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIG_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIG_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIG_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIG_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIH_PS10G_2_B_start                   : std_logic;
  signal IL_L1PHIH_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIH_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIH_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIH_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIH_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIH_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIH_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIH_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIH_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIH_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_PS10G_2_A_start                   : std_logic;
  signal IL_D2PHIA_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_PS10G_2_A_start                   : std_logic;
  signal IL_D2PHIB_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_PS10G_2_B_start                   : std_logic;
  signal IL_D2PHIB_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_PS10G_2_A_start                   : std_logic;
  signal IL_D2PHIC_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_PS10G_2_B_start                   : std_logic;
  signal IL_D2PHIC_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_PS10G_2_B_start                   : std_logic;
  signal IL_D2PHID_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIA_PS10G_2_A_start                   : std_logic;
  signal IL_D4PHIA_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIA_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIA_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIA_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIA_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIA_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIA_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIA_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIA_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIA_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_PS10G_2_A_start                   : std_logic;
  signal IL_D4PHIB_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIB_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIB_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_PS10G_2_B_start                   : std_logic;
  signal IL_D4PHIB_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIB_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIB_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_PS10G_2_A_start                   : std_logic;
  signal IL_D4PHIC_PS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_PS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_PS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIC_PS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIC_PS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_PS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_PS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_PS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_PS10G_2_B_start                   : std_logic;
  signal IL_D4PHIC_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIC_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIC_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHID_PS10G_2_B_start                   : std_logic;
  signal IL_D4PHID_PS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHID_PS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHID_PS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHID_PS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHID_PS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHID_PS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHID_PS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHID_PS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHID_PS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHID_PS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIA_PS10G_3_A_start                   : std_logic;
  signal IL_L2PHIA_PS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIA_PS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIA_PS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIA_PS10G_3_A_wea          : t_IL_36_1b;
  signal IL_L2PHIA_PS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIA_PS10G_3_A_din         : t_IL_36_DATA;
  signal IL_L2PHIA_PS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIA_PS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIA_PS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIA_PS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIB_PS10G_3_A_start                   : std_logic;
  signal IL_L2PHIB_PS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIB_PS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIB_PS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIB_PS10G_3_A_wea          : t_IL_36_1b;
  signal IL_L2PHIB_PS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIB_PS10G_3_A_din         : t_IL_36_DATA;
  signal IL_L2PHIB_PS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIB_PS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIB_PS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIB_PS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIB_PS10G_3_B_start                   : std_logic;
  signal IL_L2PHIB_PS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIB_PS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIB_PS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIB_PS10G_3_B_wea          : t_IL_36_1b;
  signal IL_L2PHIB_PS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIB_PS10G_3_B_din         : t_IL_36_DATA;
  signal IL_L2PHIB_PS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIB_PS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIB_PS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIB_PS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIC_PS10G_3_A_start                   : std_logic;
  signal IL_L2PHIC_PS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIC_PS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIC_PS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIC_PS10G_3_A_wea          : t_IL_36_1b;
  signal IL_L2PHIC_PS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIC_PS10G_3_A_din         : t_IL_36_DATA;
  signal IL_L2PHIC_PS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIC_PS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIC_PS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIC_PS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIC_PS10G_3_B_start                   : std_logic;
  signal IL_L2PHIC_PS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIC_PS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIC_PS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIC_PS10G_3_B_wea          : t_IL_36_1b;
  signal IL_L2PHIC_PS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIC_PS10G_3_B_din         : t_IL_36_DATA;
  signal IL_L2PHIC_PS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIC_PS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIC_PS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIC_PS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHID_PS10G_3_B_start                   : std_logic;
  signal IL_L2PHID_PS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L2PHID_PS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHID_PS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L2PHID_PS10G_3_B_wea          : t_IL_36_1b;
  signal IL_L2PHID_PS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHID_PS10G_3_B_din         : t_IL_36_DATA;
  signal IL_L2PHID_PS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L2PHID_PS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHID_PS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L2PHID_PS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_PS10G_3_A_start                   : std_logic;
  signal IL_D2PHIA_PS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_PS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_PS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_PS10G_3_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_PS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_PS10G_3_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_PS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_PS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_PS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_PS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_PS10G_3_A_start                   : std_logic;
  signal IL_D2PHIB_PS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_3_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_3_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_PS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_PS10G_3_B_start                   : std_logic;
  signal IL_D2PHIB_PS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_3_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_PS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_3_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_PS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_PS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_PS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_PS10G_3_A_start                   : std_logic;
  signal IL_D2PHIC_PS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_3_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_3_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_PS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_PS10G_3_B_start                   : std_logic;
  signal IL_D2PHIC_PS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_3_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_PS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_3_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_PS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_PS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_PS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_PS10G_3_B_start                   : std_logic;
  signal IL_D2PHID_PS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_PS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_PS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_PS10G_3_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_PS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_PS10G_3_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_PS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_PS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_PS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_PS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIA_PS10G_4_A_start                   : std_logic;
  signal IL_D1PHIA_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIA_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIA_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIA_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D1PHIA_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIA_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D1PHIA_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIA_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIA_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIA_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_PS10G_4_A_start                   : std_logic;
  signal IL_D1PHIB_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_PS10G_4_B_start                   : std_logic;
  signal IL_D1PHIB_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D1PHIB_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_PS10G_4_A_start                   : std_logic;
  signal IL_D1PHIC_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_PS10G_4_B_start                   : std_logic;
  signal IL_D1PHIC_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D1PHIC_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHID_PS10G_4_B_start                   : std_logic;
  signal IL_D1PHID_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHID_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHID_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHID_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D1PHID_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHID_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D1PHID_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHID_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHID_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHID_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIA_PS10G_4_A_start                   : std_logic;
  signal IL_D3PHIA_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIA_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIA_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIA_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIA_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIA_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIA_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIA_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIA_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIA_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_PS10G_4_A_start                   : std_logic;
  signal IL_D3PHIB_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_PS10G_4_B_start                   : std_logic;
  signal IL_D3PHIB_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIB_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_PS10G_4_A_start                   : std_logic;
  signal IL_D3PHIC_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_PS10G_4_B_start                   : std_logic;
  signal IL_D3PHIC_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIC_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHID_PS10G_4_B_start                   : std_logic;
  signal IL_D3PHID_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHID_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHID_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHID_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHID_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHID_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHID_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHID_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHID_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHID_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIA_PS10G_4_A_start                   : std_logic;
  signal IL_D5PHIA_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIA_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIA_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIA_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D5PHIA_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIA_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D5PHIA_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIA_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIA_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIA_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_PS10G_4_A_start                   : std_logic;
  signal IL_D5PHIB_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_PS10G_4_B_start                   : std_logic;
  signal IL_D5PHIB_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D5PHIB_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_PS10G_4_A_start                   : std_logic;
  signal IL_D5PHIC_PS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_PS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_PS10G_4_B_start                   : std_logic;
  signal IL_D5PHIC_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D5PHIC_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHID_PS10G_4_B_start                   : std_logic;
  signal IL_D5PHID_PS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHID_PS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHID_PS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHID_PS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D5PHID_PS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHID_PS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D5PHID_PS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHID_PS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHID_PS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHID_PS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIA_PS_1_A_start                   : std_logic;
  signal IL_L3PHIA_PS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIA_PS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIA_PS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIA_PS_1_A_wea          : t_IL_36_1b;
  signal IL_L3PHIA_PS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIA_PS_1_A_din         : t_IL_36_DATA;
  signal IL_L3PHIA_PS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIA_PS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIA_PS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIA_PS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIB_PS_1_A_start                   : std_logic;
  signal IL_L3PHIB_PS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIB_PS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIB_PS_1_A_wea          : t_IL_36_1b;
  signal IL_L3PHIB_PS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_1_A_din         : t_IL_36_DATA;
  signal IL_L3PHIB_PS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIB_PS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIB_PS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIC_PS_1_B_start                   : std_logic;
  signal IL_L3PHIC_PS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIC_PS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIC_PS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIC_PS_1_B_wea          : t_IL_36_1b;
  signal IL_L3PHIC_PS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIC_PS_1_B_din         : t_IL_36_DATA;
  signal IL_L3PHIC_PS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIC_PS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIC_PS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIC_PS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHID_PS_1_B_start                   : std_logic;
  signal IL_L3PHID_PS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHID_PS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHID_PS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHID_PS_1_B_wea          : t_IL_36_1b;
  signal IL_L3PHID_PS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHID_PS_1_B_din         : t_IL_36_DATA;
  signal IL_L3PHID_PS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHID_PS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHID_PS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHID_PS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_PS_1_A_start                   : std_logic;
  signal IL_D2PHIA_PS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_PS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_PS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_PS_1_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_PS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_PS_1_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_PS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_PS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_PS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_PS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_PS_1_A_start                   : std_logic;
  signal IL_D2PHIB_PS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_PS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_PS_1_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_PS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS_1_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_PS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_PS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_PS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_PS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_PS_1_B_start                   : std_logic;
  signal IL_D2PHIB_PS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_PS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_PS_1_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_PS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_PS_1_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_PS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_PS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_PS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_PS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_PS_1_A_start                   : std_logic;
  signal IL_D2PHIC_PS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_PS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_PS_1_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_PS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS_1_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_PS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_PS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_PS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_PS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_PS_1_B_start                   : std_logic;
  signal IL_D2PHIC_PS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_PS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_PS_1_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_PS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_PS_1_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_PS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_PS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_PS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_PS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_PS_1_B_start                   : std_logic;
  signal IL_D2PHID_PS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_PS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_PS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_PS_1_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_PS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_PS_1_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_PS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_PS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_PS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_PS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIA_PS_2_A_start                   : std_logic;
  signal IL_L3PHIA_PS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIA_PS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIA_PS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIA_PS_2_A_wea          : t_IL_36_1b;
  signal IL_L3PHIA_PS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIA_PS_2_A_din         : t_IL_36_DATA;
  signal IL_L3PHIA_PS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIA_PS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIA_PS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIA_PS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIB_PS_2_A_start                   : std_logic;
  signal IL_L3PHIB_PS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIB_PS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIB_PS_2_A_wea          : t_IL_36_1b;
  signal IL_L3PHIB_PS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_2_A_din         : t_IL_36_DATA;
  signal IL_L3PHIB_PS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIB_PS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIB_PS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIB_PS_2_B_start                   : std_logic;
  signal IL_L3PHIB_PS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIB_PS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIB_PS_2_B_wea          : t_IL_36_1b;
  signal IL_L3PHIB_PS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_2_B_din         : t_IL_36_DATA;
  signal IL_L3PHIB_PS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIB_PS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIB_PS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIB_PS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIC_PS_2_B_start                   : std_logic;
  signal IL_L3PHIC_PS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIC_PS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIC_PS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIC_PS_2_B_wea          : t_IL_36_1b;
  signal IL_L3PHIC_PS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIC_PS_2_B_din         : t_IL_36_DATA;
  signal IL_L3PHIC_PS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIC_PS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIC_PS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIC_PS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHID_PS_2_B_start                   : std_logic;
  signal IL_L3PHID_PS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHID_PS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHID_PS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHID_PS_2_B_wea          : t_IL_36_1b;
  signal IL_L3PHID_PS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHID_PS_2_B_din         : t_IL_36_DATA;
  signal IL_L3PHID_PS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHID_PS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHID_PS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHID_PS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIA_PS_2_A_start                   : std_logic;
  signal IL_D4PHIA_PS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIA_PS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIA_PS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIA_PS_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIA_PS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIA_PS_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIA_PS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIA_PS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIA_PS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIA_PS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_PS_2_A_start                   : std_logic;
  signal IL_D4PHIB_PS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_PS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_PS_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIB_PS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIB_PS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_PS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_PS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_PS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_PS_2_B_start                   : std_logic;
  signal IL_D4PHIB_PS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_PS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_PS_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIB_PS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_PS_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIB_PS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_PS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_PS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_PS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_PS_2_A_start                   : std_logic;
  signal IL_D4PHIC_PS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_PS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_PS_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIC_PS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIC_PS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_PS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_PS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_PS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_PS_2_B_start                   : std_logic;
  signal IL_D4PHIC_PS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_PS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_PS_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIC_PS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_PS_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIC_PS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_PS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_PS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_PS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHID_PS_2_B_start                   : std_logic;
  signal IL_D4PHID_PS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHID_PS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHID_PS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHID_PS_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHID_PS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHID_PS_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHID_PS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHID_PS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHID_PS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHID_PS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIA_negPS10G_1_A_start                   : std_logic;
  signal IL_L1PHIA_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIA_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIA_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIA_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_L1PHIA_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIA_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_L1PHIA_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIA_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIA_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIA_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIB_negPS10G_1_A_start                   : std_logic;
  signal IL_L1PHIB_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIB_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIB_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIB_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_L1PHIB_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIB_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_L1PHIB_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIB_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIB_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIB_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHID_negPS10G_1_B_start                   : std_logic;
  signal IL_L1PHID_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHID_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_L1PHID_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHID_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIE_negPS10G_1_B_start                   : std_logic;
  signal IL_L1PHIE_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIE_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_L1PHIE_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIE_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIF_negPS10G_1_B_start                   : std_logic;
  signal IL_L1PHIF_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIF_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIF_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIF_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_L1PHIF_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIF_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_L1PHIF_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIF_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIF_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIF_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIG_negPS10G_1_B_start                   : std_logic;
  signal IL_L1PHIG_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIG_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIG_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIG_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_L1PHIG_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIG_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_L1PHIG_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIG_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIG_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIG_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIA_negPS10G_1_A_start                   : std_logic;
  signal IL_D1PHIA_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIA_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIA_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIA_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D1PHIA_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIA_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D1PHIA_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIA_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIA_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIA_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_negPS10G_1_A_start                   : std_logic;
  signal IL_D1PHIB_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_negPS10G_1_B_start                   : std_logic;
  signal IL_D1PHIB_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_negPS10G_1_A_start                   : std_logic;
  signal IL_D1PHIC_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_negPS10G_1_B_start                   : std_logic;
  signal IL_D1PHIC_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHID_negPS10G_1_B_start                   : std_logic;
  signal IL_D1PHID_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHID_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHID_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHID_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D1PHID_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHID_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D1PHID_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHID_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHID_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHID_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIA_negPS10G_1_A_start                   : std_logic;
  signal IL_D3PHIA_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIA_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIA_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIA_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D3PHIA_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIA_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D3PHIA_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIA_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIA_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIA_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_negPS10G_1_A_start                   : std_logic;
  signal IL_D3PHIB_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_negPS10G_1_B_start                   : std_logic;
  signal IL_D3PHIB_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_negPS10G_1_A_start                   : std_logic;
  signal IL_D3PHIC_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_negPS10G_1_B_start                   : std_logic;
  signal IL_D3PHIC_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHID_negPS10G_1_B_start                   : std_logic;
  signal IL_D3PHID_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHID_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHID_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHID_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D3PHID_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHID_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D3PHID_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHID_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHID_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHID_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIA_negPS10G_1_A_start                   : std_logic;
  signal IL_D5PHIA_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIA_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIA_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIA_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D5PHIA_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIA_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D5PHIA_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIA_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIA_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIA_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_negPS10G_1_A_start                   : std_logic;
  signal IL_D5PHIB_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_negPS10G_1_B_start                   : std_logic;
  signal IL_D5PHIB_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_negPS10G_1_A_start                   : std_logic;
  signal IL_D5PHIC_negPS10G_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_1_A_wea          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_1_A_din         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_negPS10G_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_negPS10G_1_B_start                   : std_logic;
  signal IL_D5PHIC_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHID_negPS10G_1_B_start                   : std_logic;
  signal IL_D5PHID_negPS10G_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHID_negPS10G_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHID_negPS10G_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHID_negPS10G_1_B_wea          : t_IL_36_1b;
  signal IL_D5PHID_negPS10G_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHID_negPS10G_1_B_din         : t_IL_36_DATA;
  signal IL_D5PHID_negPS10G_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHID_negPS10G_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHID_negPS10G_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHID_negPS10G_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIA_negPS10G_2_A_start                   : std_logic;
  signal IL_L1PHIA_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIA_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIA_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIA_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIA_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIA_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIA_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIA_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIA_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIA_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIB_negPS10G_2_A_start                   : std_logic;
  signal IL_L1PHIB_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIB_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIB_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIB_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIB_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIB_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIB_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIB_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIB_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIB_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIC_negPS10G_2_A_start                   : std_logic;
  signal IL_L1PHIC_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIC_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIC_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIC_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIC_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIC_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIC_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIC_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIC_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIC_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHID_negPS10G_2_A_start                   : std_logic;
  signal IL_L1PHID_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHID_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHID_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHID_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHID_negPS10G_2_B_start                   : std_logic;
  signal IL_L1PHID_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHID_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHID_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHID_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHID_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHID_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIE_negPS10G_2_A_start                   : std_logic;
  signal IL_L1PHIE_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIE_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_L1PHIE_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIE_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIE_negPS10G_2_B_start                   : std_logic;
  signal IL_L1PHIE_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIE_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIE_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIE_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIE_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIE_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIF_negPS10G_2_B_start                   : std_logic;
  signal IL_L1PHIF_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIF_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIF_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIF_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIF_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIF_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIF_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIF_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIF_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIF_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIG_negPS10G_2_B_start                   : std_logic;
  signal IL_L1PHIG_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIG_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIG_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIG_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIG_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIG_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIG_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIG_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIG_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIG_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L1PHIH_negPS10G_2_B_start                   : std_logic;
  signal IL_L1PHIH_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L1PHIH_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L1PHIH_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L1PHIH_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_L1PHIH_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L1PHIH_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_L1PHIH_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L1PHIH_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L1PHIH_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L1PHIH_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_negPS10G_2_A_start                   : std_logic;
  signal IL_D2PHIA_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_negPS10G_2_A_start                   : std_logic;
  signal IL_D2PHIB_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_negPS10G_2_B_start                   : std_logic;
  signal IL_D2PHIB_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_negPS10G_2_A_start                   : std_logic;
  signal IL_D2PHIC_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_negPS10G_2_B_start                   : std_logic;
  signal IL_D2PHIC_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_negPS10G_2_B_start                   : std_logic;
  signal IL_D2PHID_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIA_negPS10G_2_A_start                   : std_logic;
  signal IL_D4PHIA_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIA_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIA_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIA_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIA_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIA_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIA_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIA_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIA_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIA_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_negPS10G_2_A_start                   : std_logic;
  signal IL_D4PHIB_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIB_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_negPS10G_2_B_start                   : std_logic;
  signal IL_D4PHIB_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIB_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_negPS10G_2_A_start                   : std_logic;
  signal IL_D4PHIC_negPS10G_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_negPS10G_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS10G_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS10G_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIC_negPS10G_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS10G_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS10G_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_negPS10G_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS10G_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_negPS10G_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_negPS10G_2_B_start                   : std_logic;
  signal IL_D4PHIC_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIC_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHID_negPS10G_2_B_start                   : std_logic;
  signal IL_D4PHID_negPS10G_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHID_negPS10G_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHID_negPS10G_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHID_negPS10G_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHID_negPS10G_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHID_negPS10G_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHID_negPS10G_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHID_negPS10G_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHID_negPS10G_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHID_negPS10G_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIA_negPS10G_3_A_start                   : std_logic;
  signal IL_L2PHIA_negPS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIA_negPS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIA_negPS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIA_negPS10G_3_A_wea          : t_IL_36_1b;
  signal IL_L2PHIA_negPS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIA_negPS10G_3_A_din         : t_IL_36_DATA;
  signal IL_L2PHIA_negPS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIA_negPS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIA_negPS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIA_negPS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIB_negPS10G_3_A_start                   : std_logic;
  signal IL_L2PHIB_negPS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIB_negPS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIB_negPS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIB_negPS10G_3_A_wea          : t_IL_36_1b;
  signal IL_L2PHIB_negPS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIB_negPS10G_3_A_din         : t_IL_36_DATA;
  signal IL_L2PHIB_negPS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIB_negPS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIB_negPS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIB_negPS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIB_negPS10G_3_B_start                   : std_logic;
  signal IL_L2PHIB_negPS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIB_negPS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIB_negPS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIB_negPS10G_3_B_wea          : t_IL_36_1b;
  signal IL_L2PHIB_negPS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIB_negPS10G_3_B_din         : t_IL_36_DATA;
  signal IL_L2PHIB_negPS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIB_negPS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIB_negPS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIB_negPS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIC_negPS10G_3_A_start                   : std_logic;
  signal IL_L2PHIC_negPS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIC_negPS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIC_negPS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIC_negPS10G_3_A_wea          : t_IL_36_1b;
  signal IL_L2PHIC_negPS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIC_negPS10G_3_A_din         : t_IL_36_DATA;
  signal IL_L2PHIC_negPS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIC_negPS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIC_negPS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIC_negPS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHIC_negPS10G_3_B_start                   : std_logic;
  signal IL_L2PHIC_negPS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L2PHIC_negPS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHIC_negPS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L2PHIC_negPS10G_3_B_wea          : t_IL_36_1b;
  signal IL_L2PHIC_negPS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHIC_negPS10G_3_B_din         : t_IL_36_DATA;
  signal IL_L2PHIC_negPS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L2PHIC_negPS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHIC_negPS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L2PHIC_negPS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L2PHID_negPS10G_3_B_start                   : std_logic;
  signal IL_L2PHID_negPS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L2PHID_negPS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L2PHID_negPS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L2PHID_negPS10G_3_B_wea          : t_IL_36_1b;
  signal IL_L2PHID_negPS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L2PHID_negPS10G_3_B_din         : t_IL_36_DATA;
  signal IL_L2PHID_negPS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L2PHID_negPS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L2PHID_negPS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L2PHID_negPS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_negPS10G_3_A_start                   : std_logic;
  signal IL_D2PHIA_negPS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_negPS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_negPS10G_3_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_negPS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS10G_3_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_negPS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_negPS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_negPS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_negPS10G_3_A_start                   : std_logic;
  signal IL_D2PHIB_negPS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_3_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_3_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_negPS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_negPS10G_3_B_start                   : std_logic;
  signal IL_D2PHIB_negPS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_3_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_negPS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_3_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_negPS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_negPS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_negPS10G_3_A_start                   : std_logic;
  signal IL_D2PHIC_negPS10G_3_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_3_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_3_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_3_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_3_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_negPS10G_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_3_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_negPS10G_3_B_start                   : std_logic;
  signal IL_D2PHIC_negPS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_3_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_negPS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_3_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_negPS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_negPS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_negPS10G_3_B_start                   : std_logic;
  signal IL_D2PHID_negPS10G_3_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_negPS10G_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_negPS10G_3_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_negPS10G_3_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_negPS10G_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_negPS10G_3_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_negPS10G_3_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_negPS10G_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_negPS10G_3_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_negPS10G_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIA_negPS10G_4_A_start                   : std_logic;
  signal IL_D1PHIA_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIA_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIA_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIA_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D1PHIA_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIA_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D1PHIA_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIA_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIA_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIA_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_negPS10G_4_A_start                   : std_logic;
  signal IL_D1PHIB_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_negPS10G_4_B_start                   : std_logic;
  signal IL_D1PHIB_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D1PHIB_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_negPS10G_4_A_start                   : std_logic;
  signal IL_D1PHIC_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_negPS10G_4_B_start                   : std_logic;
  signal IL_D1PHIC_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D1PHIC_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHID_negPS10G_4_B_start                   : std_logic;
  signal IL_D1PHID_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHID_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHID_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHID_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D1PHID_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHID_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D1PHID_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHID_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHID_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHID_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIA_negPS10G_4_A_start                   : std_logic;
  signal IL_D3PHIA_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIA_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIA_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIA_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIA_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIA_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIA_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIA_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIA_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIA_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_negPS10G_4_A_start                   : std_logic;
  signal IL_D3PHIB_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_negPS10G_4_B_start                   : std_logic;
  signal IL_D3PHIB_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIB_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_negPS10G_4_A_start                   : std_logic;
  signal IL_D3PHIC_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_negPS10G_4_B_start                   : std_logic;
  signal IL_D3PHIC_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIC_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHID_negPS10G_4_B_start                   : std_logic;
  signal IL_D3PHID_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHID_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHID_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHID_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHID_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHID_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHID_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHID_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHID_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHID_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIA_negPS10G_4_A_start                   : std_logic;
  signal IL_D5PHIA_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIA_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIA_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIA_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D5PHIA_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIA_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D5PHIA_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIA_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIA_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIA_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_negPS10G_4_A_start                   : std_logic;
  signal IL_D5PHIB_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_negPS10G_4_B_start                   : std_logic;
  signal IL_D5PHIB_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D5PHIB_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_negPS10G_4_A_start                   : std_logic;
  signal IL_D5PHIC_negPS10G_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_4_A_wea          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_4_A_din         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_negPS10G_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_negPS10G_4_B_start                   : std_logic;
  signal IL_D5PHIC_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D5PHIC_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHID_negPS10G_4_B_start                   : std_logic;
  signal IL_D5PHID_negPS10G_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHID_negPS10G_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHID_negPS10G_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHID_negPS10G_4_B_wea          : t_IL_36_1b;
  signal IL_D5PHID_negPS10G_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHID_negPS10G_4_B_din         : t_IL_36_DATA;
  signal IL_D5PHID_negPS10G_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHID_negPS10G_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHID_negPS10G_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHID_negPS10G_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIA_negPS_1_A_start                   : std_logic;
  signal IL_L3PHIA_negPS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIA_negPS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIA_negPS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIA_negPS_1_A_wea          : t_IL_36_1b;
  signal IL_L3PHIA_negPS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIA_negPS_1_A_din         : t_IL_36_DATA;
  signal IL_L3PHIA_negPS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIA_negPS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIA_negPS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIA_negPS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIB_negPS_1_A_start                   : std_logic;
  signal IL_L3PHIB_negPS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_1_A_wea          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_1_A_din         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIB_negPS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIB_negPS_1_B_start                   : std_logic;
  signal IL_L3PHIB_negPS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_1_B_wea          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_1_B_din         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIB_negPS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIC_negPS_1_B_start                   : std_logic;
  signal IL_L3PHIC_negPS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIC_negPS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIC_negPS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIC_negPS_1_B_wea          : t_IL_36_1b;
  signal IL_L3PHIC_negPS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIC_negPS_1_B_din         : t_IL_36_DATA;
  signal IL_L3PHIC_negPS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIC_negPS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIC_negPS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIC_negPS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHID_negPS_1_B_start                   : std_logic;
  signal IL_L3PHID_negPS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHID_negPS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHID_negPS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHID_negPS_1_B_wea          : t_IL_36_1b;
  signal IL_L3PHID_negPS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHID_negPS_1_B_din         : t_IL_36_DATA;
  signal IL_L3PHID_negPS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHID_negPS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHID_negPS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHID_negPS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_negPS_1_A_start                   : std_logic;
  signal IL_D2PHIA_negPS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_negPS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_negPS_1_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_negPS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS_1_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_negPS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_negPS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_negPS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_negPS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_negPS_1_A_start                   : std_logic;
  signal IL_D2PHIB_negPS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_negPS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS_1_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_negPS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS_1_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_negPS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_negPS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_negPS_1_B_start                   : std_logic;
  signal IL_D2PHIB_negPS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_negPS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS_1_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_negPS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS_1_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_negPS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_negPS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_negPS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_negPS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_negPS_1_A_start                   : std_logic;
  signal IL_D2PHIC_negPS_1_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_negPS_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS_1_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS_1_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_negPS_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS_1_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS_1_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_negPS_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS_1_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_negPS_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_negPS_1_B_start                   : std_logic;
  signal IL_D2PHIC_negPS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_negPS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS_1_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_negPS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS_1_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_negPS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_negPS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_negPS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_negPS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_negPS_1_B_start                   : std_logic;
  signal IL_D2PHID_negPS_1_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_negPS_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_negPS_1_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_negPS_1_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_negPS_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_negPS_1_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_negPS_1_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_negPS_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_negPS_1_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_negPS_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIA_negPS_2_A_start                   : std_logic;
  signal IL_L3PHIA_negPS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIA_negPS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIA_negPS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIA_negPS_2_A_wea          : t_IL_36_1b;
  signal IL_L3PHIA_negPS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIA_negPS_2_A_din         : t_IL_36_DATA;
  signal IL_L3PHIA_negPS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIA_negPS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIA_negPS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIA_negPS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIB_negPS_2_A_start                   : std_logic;
  signal IL_L3PHIB_negPS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_2_A_wea          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_2_A_din         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIB_negPS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIB_negPS_2_B_start                   : std_logic;
  signal IL_L3PHIB_negPS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_2_B_wea          : t_IL_36_1b;
  signal IL_L3PHIB_negPS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_2_B_din         : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIB_negPS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIB_negPS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIB_negPS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHIC_negPS_2_B_start                   : std_logic;
  signal IL_L3PHIC_negPS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHIC_negPS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHIC_negPS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHIC_negPS_2_B_wea          : t_IL_36_1b;
  signal IL_L3PHIC_negPS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHIC_negPS_2_B_din         : t_IL_36_DATA;
  signal IL_L3PHIC_negPS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHIC_negPS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHIC_negPS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHIC_negPS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L3PHID_negPS_2_B_start                   : std_logic;
  signal IL_L3PHID_negPS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L3PHID_negPS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L3PHID_negPS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L3PHID_negPS_2_B_wea          : t_IL_36_1b;
  signal IL_L3PHID_negPS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L3PHID_negPS_2_B_din         : t_IL_36_DATA;
  signal IL_L3PHID_negPS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L3PHID_negPS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L3PHID_negPS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L3PHID_negPS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIA_negPS_2_A_start                   : std_logic;
  signal IL_D4PHIA_negPS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIA_negPS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIA_negPS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIA_negPS_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIA_negPS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIA_negPS_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIA_negPS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIA_negPS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIA_negPS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIA_negPS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_negPS_2_A_start                   : std_logic;
  signal IL_D4PHIB_negPS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_negPS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIB_negPS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_negPS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_negPS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_negPS_2_B_start                   : std_logic;
  signal IL_D4PHIB_negPS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_negPS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIB_negPS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIB_negPS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_negPS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_negPS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_negPS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_negPS_2_A_start                   : std_logic;
  signal IL_D4PHIC_negPS_2_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_negPS_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS_2_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS_2_A_wea          : t_IL_36_1b;
  signal IL_D4PHIC_negPS_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS_2_A_din         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS_2_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_negPS_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS_2_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_negPS_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_negPS_2_B_start                   : std_logic;
  signal IL_D4PHIC_negPS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_negPS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHIC_negPS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHIC_negPS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_negPS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_negPS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_negPS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHID_negPS_2_B_start                   : std_logic;
  signal IL_D4PHID_negPS_2_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHID_negPS_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHID_negPS_2_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHID_negPS_2_B_wea          : t_IL_36_1b;
  signal IL_D4PHID_negPS_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHID_negPS_2_B_din         : t_IL_36_DATA;
  signal IL_D4PHID_negPS_2_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHID_negPS_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHID_negPS_2_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHID_negPS_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIA_2S_1_A_start                   : std_logic;
  signal IL_L4PHIA_2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIA_2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIA_2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIA_2S_1_A_wea          : t_IL_36_1b;
  signal IL_L4PHIA_2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIA_2S_1_A_din         : t_IL_36_DATA;
  signal IL_L4PHIA_2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIA_2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIA_2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIA_2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIB_2S_1_A_start                   : std_logic;
  signal IL_L4PHIB_2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIB_2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIB_2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIB_2S_1_A_wea          : t_IL_36_1b;
  signal IL_L4PHIB_2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIB_2S_1_A_din         : t_IL_36_DATA;
  signal IL_L4PHIB_2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIB_2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIB_2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIB_2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIB_2S_1_B_start                   : std_logic;
  signal IL_L4PHIB_2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIB_2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIB_2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIB_2S_1_B_wea          : t_IL_36_1b;
  signal IL_L4PHIB_2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIB_2S_1_B_din         : t_IL_36_DATA;
  signal IL_L4PHIB_2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIB_2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIB_2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIB_2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIC_2S_1_A_start                   : std_logic;
  signal IL_L4PHIC_2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIC_2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIC_2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIC_2S_1_A_wea          : t_IL_36_1b;
  signal IL_L4PHIC_2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIC_2S_1_A_din         : t_IL_36_DATA;
  signal IL_L4PHIC_2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIC_2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIC_2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIC_2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIC_2S_1_B_start                   : std_logic;
  signal IL_L4PHIC_2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIC_2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIC_2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIC_2S_1_B_wea          : t_IL_36_1b;
  signal IL_L4PHIC_2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIC_2S_1_B_din         : t_IL_36_DATA;
  signal IL_L4PHIC_2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIC_2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIC_2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIC_2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHID_2S_1_B_start                   : std_logic;
  signal IL_L4PHID_2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L4PHID_2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHID_2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L4PHID_2S_1_B_wea          : t_IL_36_1b;
  signal IL_L4PHID_2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHID_2S_1_B_din         : t_IL_36_DATA;
  signal IL_L4PHID_2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L4PHID_2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHID_2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L4PHID_2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIA_2S_1_A_start                   : std_logic;
  signal IL_L5PHIA_2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIA_2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIA_2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIA_2S_1_A_wea          : t_IL_36_1b;
  signal IL_L5PHIA_2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIA_2S_1_A_din         : t_IL_36_DATA;
  signal IL_L5PHIA_2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIA_2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIA_2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIA_2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHID_2S_1_B_start                   : std_logic;
  signal IL_L5PHID_2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHID_2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHID_2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHID_2S_1_B_wea          : t_IL_36_1b;
  signal IL_L5PHID_2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHID_2S_1_B_din         : t_IL_36_DATA;
  signal IL_L5PHID_2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHID_2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHID_2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHID_2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIA_2S_2_A_start                   : std_logic;
  signal IL_L5PHIA_2S_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIA_2S_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIA_2S_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIA_2S_2_A_wea          : t_IL_36_1b;
  signal IL_L5PHIA_2S_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIA_2S_2_A_din         : t_IL_36_DATA;
  signal IL_L5PHIA_2S_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIA_2S_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIA_2S_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIA_2S_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIB_2S_2_A_start                   : std_logic;
  signal IL_L5PHIB_2S_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIB_2S_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIB_2S_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIB_2S_2_A_wea          : t_IL_36_1b;
  signal IL_L5PHIB_2S_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIB_2S_2_A_din         : t_IL_36_DATA;
  signal IL_L5PHIB_2S_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIB_2S_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIB_2S_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIB_2S_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIB_2S_2_B_start                   : std_logic;
  signal IL_L5PHIB_2S_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIB_2S_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIB_2S_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIB_2S_2_B_wea          : t_IL_36_1b;
  signal IL_L5PHIB_2S_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIB_2S_2_B_din         : t_IL_36_DATA;
  signal IL_L5PHIB_2S_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIB_2S_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIB_2S_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIB_2S_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIC_2S_2_A_start                   : std_logic;
  signal IL_L5PHIC_2S_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIC_2S_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIC_2S_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIC_2S_2_A_wea          : t_IL_36_1b;
  signal IL_L5PHIC_2S_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIC_2S_2_A_din         : t_IL_36_DATA;
  signal IL_L5PHIC_2S_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIC_2S_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIC_2S_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIC_2S_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIC_2S_2_B_start                   : std_logic;
  signal IL_L5PHIC_2S_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIC_2S_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIC_2S_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIC_2S_2_B_wea          : t_IL_36_1b;
  signal IL_L5PHIC_2S_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIC_2S_2_B_din         : t_IL_36_DATA;
  signal IL_L5PHIC_2S_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIC_2S_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIC_2S_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIC_2S_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHID_2S_2_B_start                   : std_logic;
  signal IL_L5PHID_2S_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHID_2S_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHID_2S_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHID_2S_2_B_wea          : t_IL_36_1b;
  signal IL_L5PHID_2S_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHID_2S_2_B_din         : t_IL_36_DATA;
  signal IL_L5PHID_2S_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHID_2S_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHID_2S_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHID_2S_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIA_2S_3_A_start                   : std_logic;
  signal IL_L6PHIA_2S_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIA_2S_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIA_2S_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIA_2S_3_A_wea          : t_IL_36_1b;
  signal IL_L6PHIA_2S_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIA_2S_3_A_din         : t_IL_36_DATA;
  signal IL_L6PHIA_2S_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIA_2S_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIA_2S_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIA_2S_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIB_2S_3_A_start                   : std_logic;
  signal IL_L6PHIB_2S_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIB_2S_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIB_2S_3_A_wea          : t_IL_36_1b;
  signal IL_L6PHIB_2S_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_3_A_din         : t_IL_36_DATA;
  signal IL_L6PHIB_2S_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIB_2S_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIB_2S_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIC_2S_3_A_start                   : std_logic;
  signal IL_L6PHIC_2S_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIC_2S_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIC_2S_3_A_wea          : t_IL_36_1b;
  signal IL_L6PHIC_2S_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_3_A_din         : t_IL_36_DATA;
  signal IL_L6PHIC_2S_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIC_2S_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIC_2S_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIC_2S_3_B_start                   : std_logic;
  signal IL_L6PHIC_2S_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIC_2S_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIC_2S_3_B_wea          : t_IL_36_1b;
  signal IL_L6PHIC_2S_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_3_B_din         : t_IL_36_DATA;
  signal IL_L6PHIC_2S_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIC_2S_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIC_2S_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHID_2S_3_B_start                   : std_logic;
  signal IL_L6PHID_2S_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHID_2S_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHID_2S_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHID_2S_3_B_wea          : t_IL_36_1b;
  signal IL_L6PHID_2S_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHID_2S_3_B_din         : t_IL_36_DATA;
  signal IL_L6PHID_2S_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHID_2S_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHID_2S_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHID_2S_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIA_2S_4_A_start                   : std_logic;
  signal IL_L6PHIA_2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIA_2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIA_2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIA_2S_4_A_wea          : t_IL_36_1b;
  signal IL_L6PHIA_2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIA_2S_4_A_din         : t_IL_36_DATA;
  signal IL_L6PHIA_2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIA_2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIA_2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIA_2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIB_2S_4_A_start                   : std_logic;
  signal IL_L6PHIB_2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIB_2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIB_2S_4_A_wea          : t_IL_36_1b;
  signal IL_L6PHIB_2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_4_A_din         : t_IL_36_DATA;
  signal IL_L6PHIB_2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIB_2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIB_2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIB_2S_4_B_start                   : std_logic;
  signal IL_L6PHIB_2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIB_2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIB_2S_4_B_wea          : t_IL_36_1b;
  signal IL_L6PHIB_2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_4_B_din         : t_IL_36_DATA;
  signal IL_L6PHIB_2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIB_2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIB_2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIB_2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIC_2S_4_B_start                   : std_logic;
  signal IL_L6PHIC_2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIC_2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIC_2S_4_B_wea          : t_IL_36_1b;
  signal IL_L6PHIC_2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_4_B_din         : t_IL_36_DATA;
  signal IL_L6PHIC_2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIC_2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIC_2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIC_2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHID_2S_4_B_start                   : std_logic;
  signal IL_L6PHID_2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHID_2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHID_2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHID_2S_4_B_wea          : t_IL_36_1b;
  signal IL_L6PHID_2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHID_2S_4_B_din         : t_IL_36_DATA;
  signal IL_L6PHID_2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHID_2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHID_2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHID_2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIA_2S_4_A_start                   : std_logic;
  signal IL_D3PHIA_2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIA_2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIA_2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIA_2S_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIA_2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIA_2S_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIA_2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIA_2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIA_2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIA_2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_2S_4_A_start                   : std_logic;
  signal IL_D3PHIB_2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_2S_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIB_2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_2S_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIB_2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_2S_4_B_start                   : std_logic;
  signal IL_D3PHIB_2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_2S_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIB_2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_2S_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIB_2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_2S_4_A_start                   : std_logic;
  signal IL_D3PHIC_2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_2S_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIC_2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_2S_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIC_2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_2S_4_B_start                   : std_logic;
  signal IL_D3PHIC_2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_2S_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIC_2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_2S_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIC_2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHID_2S_4_B_start                   : std_logic;
  signal IL_D3PHID_2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHID_2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHID_2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHID_2S_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHID_2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHID_2S_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHID_2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHID_2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHID_2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHID_2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIA_2S_5_A_start                   : std_logic;
  signal IL_D1PHIA_2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIA_2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIA_2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIA_2S_5_A_wea          : t_IL_36_1b;
  signal IL_D1PHIA_2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIA_2S_5_A_din         : t_IL_36_DATA;
  signal IL_D1PHIA_2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIA_2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIA_2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIA_2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_2S_5_A_start                   : std_logic;
  signal IL_D1PHIB_2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_2S_5_A_wea          : t_IL_36_1b;
  signal IL_D1PHIB_2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_2S_5_A_din         : t_IL_36_DATA;
  signal IL_D1PHIB_2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_2S_5_B_start                   : std_logic;
  signal IL_D1PHIB_2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_2S_5_B_wea          : t_IL_36_1b;
  signal IL_D1PHIB_2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_2S_5_B_din         : t_IL_36_DATA;
  signal IL_D1PHIB_2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_2S_5_A_start                   : std_logic;
  signal IL_D1PHIC_2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_2S_5_A_wea          : t_IL_36_1b;
  signal IL_D1PHIC_2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_2S_5_A_din         : t_IL_36_DATA;
  signal IL_D1PHIC_2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_2S_5_B_start                   : std_logic;
  signal IL_D1PHIC_2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_2S_5_B_wea          : t_IL_36_1b;
  signal IL_D1PHIC_2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_2S_5_B_din         : t_IL_36_DATA;
  signal IL_D1PHIC_2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHID_2S_5_B_start                   : std_logic;
  signal IL_D1PHID_2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHID_2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHID_2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHID_2S_5_B_wea          : t_IL_36_1b;
  signal IL_D1PHID_2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHID_2S_5_B_din         : t_IL_36_DATA;
  signal IL_D1PHID_2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHID_2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHID_2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHID_2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIA_2S_5_A_start                   : std_logic;
  signal IL_D4PHIA_2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIA_2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIA_2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIA_2S_5_A_wea          : t_IL_36_1b;
  signal IL_D4PHIA_2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIA_2S_5_A_din         : t_IL_36_DATA;
  signal IL_D4PHIA_2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIA_2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIA_2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIA_2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_2S_5_A_start                   : std_logic;
  signal IL_D4PHIB_2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_2S_5_A_wea          : t_IL_36_1b;
  signal IL_D4PHIB_2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_2S_5_A_din         : t_IL_36_DATA;
  signal IL_D4PHIB_2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_2S_5_B_start                   : std_logic;
  signal IL_D4PHIB_2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_2S_5_B_wea          : t_IL_36_1b;
  signal IL_D4PHIB_2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_2S_5_B_din         : t_IL_36_DATA;
  signal IL_D4PHIB_2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_2S_5_A_start                   : std_logic;
  signal IL_D4PHIC_2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_2S_5_A_wea          : t_IL_36_1b;
  signal IL_D4PHIC_2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_2S_5_A_din         : t_IL_36_DATA;
  signal IL_D4PHIC_2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_2S_5_B_start                   : std_logic;
  signal IL_D4PHIC_2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_2S_5_B_wea          : t_IL_36_1b;
  signal IL_D4PHIC_2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_2S_5_B_din         : t_IL_36_DATA;
  signal IL_D4PHIC_2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHID_2S_5_B_start                   : std_logic;
  signal IL_D4PHID_2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHID_2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHID_2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHID_2S_5_B_wea          : t_IL_36_1b;
  signal IL_D4PHID_2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHID_2S_5_B_din         : t_IL_36_DATA;
  signal IL_D4PHID_2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHID_2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHID_2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHID_2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_2S_6_A_start                   : std_logic;
  signal IL_D2PHIA_2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_2S_6_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_2S_6_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_2S_6_A_start                   : std_logic;
  signal IL_D2PHIB_2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_2S_6_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_2S_6_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_2S_6_B_start                   : std_logic;
  signal IL_D2PHIB_2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_2S_6_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_2S_6_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_2S_6_A_start                   : std_logic;
  signal IL_D2PHIC_2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_2S_6_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_2S_6_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_2S_6_B_start                   : std_logic;
  signal IL_D2PHIC_2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_2S_6_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_2S_6_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_2S_6_B_start                   : std_logic;
  signal IL_D2PHID_2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_2S_6_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_2S_6_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIA_2S_6_A_start                   : std_logic;
  signal IL_D5PHIA_2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIA_2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIA_2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIA_2S_6_A_wea          : t_IL_36_1b;
  signal IL_D5PHIA_2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIA_2S_6_A_din         : t_IL_36_DATA;
  signal IL_D5PHIA_2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIA_2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIA_2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIA_2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_2S_6_A_start                   : std_logic;
  signal IL_D5PHIB_2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_2S_6_A_wea          : t_IL_36_1b;
  signal IL_D5PHIB_2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_2S_6_A_din         : t_IL_36_DATA;
  signal IL_D5PHIB_2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_2S_6_B_start                   : std_logic;
  signal IL_D5PHIB_2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_2S_6_B_wea          : t_IL_36_1b;
  signal IL_D5PHIB_2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_2S_6_B_din         : t_IL_36_DATA;
  signal IL_D5PHIB_2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_2S_6_A_start                   : std_logic;
  signal IL_D5PHIC_2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_2S_6_A_wea          : t_IL_36_1b;
  signal IL_D5PHIC_2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_2S_6_A_din         : t_IL_36_DATA;
  signal IL_D5PHIC_2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_2S_6_B_start                   : std_logic;
  signal IL_D5PHIC_2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_2S_6_B_wea          : t_IL_36_1b;
  signal IL_D5PHIC_2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_2S_6_B_din         : t_IL_36_DATA;
  signal IL_D5PHIC_2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHID_2S_6_B_start                   : std_logic;
  signal IL_D5PHID_2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHID_2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHID_2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHID_2S_6_B_wea          : t_IL_36_1b;
  signal IL_D5PHID_2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHID_2S_6_B_din         : t_IL_36_DATA;
  signal IL_D5PHID_2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHID_2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHID_2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHID_2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIA_neg2S_1_A_start                   : std_logic;
  signal IL_L4PHIA_neg2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIA_neg2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIA_neg2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIA_neg2S_1_A_wea          : t_IL_36_1b;
  signal IL_L4PHIA_neg2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIA_neg2S_1_A_din         : t_IL_36_DATA;
  signal IL_L4PHIA_neg2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIA_neg2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIA_neg2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIA_neg2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIB_neg2S_1_A_start                   : std_logic;
  signal IL_L4PHIB_neg2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIB_neg2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIB_neg2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIB_neg2S_1_A_wea          : t_IL_36_1b;
  signal IL_L4PHIB_neg2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIB_neg2S_1_A_din         : t_IL_36_DATA;
  signal IL_L4PHIB_neg2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIB_neg2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIB_neg2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIB_neg2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIB_neg2S_1_B_start                   : std_logic;
  signal IL_L4PHIB_neg2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIB_neg2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIB_neg2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIB_neg2S_1_B_wea          : t_IL_36_1b;
  signal IL_L4PHIB_neg2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIB_neg2S_1_B_din         : t_IL_36_DATA;
  signal IL_L4PHIB_neg2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIB_neg2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIB_neg2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIB_neg2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIC_neg2S_1_A_start                   : std_logic;
  signal IL_L4PHIC_neg2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIC_neg2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIC_neg2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIC_neg2S_1_A_wea          : t_IL_36_1b;
  signal IL_L4PHIC_neg2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIC_neg2S_1_A_din         : t_IL_36_DATA;
  signal IL_L4PHIC_neg2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIC_neg2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIC_neg2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIC_neg2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHIC_neg2S_1_B_start                   : std_logic;
  signal IL_L4PHIC_neg2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L4PHIC_neg2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHIC_neg2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L4PHIC_neg2S_1_B_wea          : t_IL_36_1b;
  signal IL_L4PHIC_neg2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHIC_neg2S_1_B_din         : t_IL_36_DATA;
  signal IL_L4PHIC_neg2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L4PHIC_neg2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHIC_neg2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L4PHIC_neg2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L4PHID_neg2S_1_B_start                   : std_logic;
  signal IL_L4PHID_neg2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L4PHID_neg2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L4PHID_neg2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L4PHID_neg2S_1_B_wea          : t_IL_36_1b;
  signal IL_L4PHID_neg2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L4PHID_neg2S_1_B_din         : t_IL_36_DATA;
  signal IL_L4PHID_neg2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L4PHID_neg2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L4PHID_neg2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L4PHID_neg2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIA_neg2S_1_A_start                   : std_logic;
  signal IL_L5PHIA_neg2S_1_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIA_neg2S_1_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIA_neg2S_1_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIA_neg2S_1_A_wea          : t_IL_36_1b;
  signal IL_L5PHIA_neg2S_1_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIA_neg2S_1_A_din         : t_IL_36_DATA;
  signal IL_L5PHIA_neg2S_1_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIA_neg2S_1_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIA_neg2S_1_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIA_neg2S_1_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHID_neg2S_1_B_start                   : std_logic;
  signal IL_L5PHID_neg2S_1_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHID_neg2S_1_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHID_neg2S_1_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHID_neg2S_1_B_wea          : t_IL_36_1b;
  signal IL_L5PHID_neg2S_1_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHID_neg2S_1_B_din         : t_IL_36_DATA;
  signal IL_L5PHID_neg2S_1_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHID_neg2S_1_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHID_neg2S_1_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHID_neg2S_1_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIA_neg2S_2_A_start                   : std_logic;
  signal IL_L5PHIA_neg2S_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIA_neg2S_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIA_neg2S_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIA_neg2S_2_A_wea          : t_IL_36_1b;
  signal IL_L5PHIA_neg2S_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIA_neg2S_2_A_din         : t_IL_36_DATA;
  signal IL_L5PHIA_neg2S_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIA_neg2S_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIA_neg2S_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIA_neg2S_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIB_neg2S_2_A_start                   : std_logic;
  signal IL_L5PHIB_neg2S_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIB_neg2S_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIB_neg2S_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIB_neg2S_2_A_wea          : t_IL_36_1b;
  signal IL_L5PHIB_neg2S_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIB_neg2S_2_A_din         : t_IL_36_DATA;
  signal IL_L5PHIB_neg2S_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIB_neg2S_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIB_neg2S_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIB_neg2S_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIB_neg2S_2_B_start                   : std_logic;
  signal IL_L5PHIB_neg2S_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIB_neg2S_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIB_neg2S_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIB_neg2S_2_B_wea          : t_IL_36_1b;
  signal IL_L5PHIB_neg2S_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIB_neg2S_2_B_din         : t_IL_36_DATA;
  signal IL_L5PHIB_neg2S_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIB_neg2S_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIB_neg2S_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIB_neg2S_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIC_neg2S_2_A_start                   : std_logic;
  signal IL_L5PHIC_neg2S_2_A_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIC_neg2S_2_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIC_neg2S_2_A_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIC_neg2S_2_A_wea          : t_IL_36_1b;
  signal IL_L5PHIC_neg2S_2_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIC_neg2S_2_A_din         : t_IL_36_DATA;
  signal IL_L5PHIC_neg2S_2_A_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIC_neg2S_2_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIC_neg2S_2_A_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIC_neg2S_2_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHIC_neg2S_2_B_start                   : std_logic;
  signal IL_L5PHIC_neg2S_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHIC_neg2S_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHIC_neg2S_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHIC_neg2S_2_B_wea          : t_IL_36_1b;
  signal IL_L5PHIC_neg2S_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHIC_neg2S_2_B_din         : t_IL_36_DATA;
  signal IL_L5PHIC_neg2S_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHIC_neg2S_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHIC_neg2S_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHIC_neg2S_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L5PHID_neg2S_2_B_start                   : std_logic;
  signal IL_L5PHID_neg2S_2_B_wea_delay          : t_IL_36_1b;
  signal IL_L5PHID_neg2S_2_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L5PHID_neg2S_2_B_din_delay         : t_IL_36_DATA;
  signal IL_L5PHID_neg2S_2_B_wea          : t_IL_36_1b;
  signal IL_L5PHID_neg2S_2_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L5PHID_neg2S_2_B_din         : t_IL_36_DATA;
  signal IL_L5PHID_neg2S_2_B_enb          : t_IL_36_1b := '1';
  signal IL_L5PHID_neg2S_2_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L5PHID_neg2S_2_B_V_dout        : t_IL_36_DATA;
  signal IL_L5PHID_neg2S_2_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIA_neg2S_3_A_start                   : std_logic;
  signal IL_L6PHIA_neg2S_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIA_neg2S_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIA_neg2S_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIA_neg2S_3_A_wea          : t_IL_36_1b;
  signal IL_L6PHIA_neg2S_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIA_neg2S_3_A_din         : t_IL_36_DATA;
  signal IL_L6PHIA_neg2S_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIA_neg2S_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIA_neg2S_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIA_neg2S_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIB_neg2S_3_A_start                   : std_logic;
  signal IL_L6PHIB_neg2S_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIB_neg2S_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_3_A_wea          : t_IL_36_1b;
  signal IL_L6PHIB_neg2S_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_3_A_din         : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIB_neg2S_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIC_neg2S_3_A_start                   : std_logic;
  signal IL_L6PHIC_neg2S_3_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIC_neg2S_3_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_3_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_3_A_wea          : t_IL_36_1b;
  signal IL_L6PHIC_neg2S_3_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_3_A_din         : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_3_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIC_neg2S_3_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_3_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_3_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIC_neg2S_3_B_start                   : std_logic;
  signal IL_L6PHIC_neg2S_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIC_neg2S_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_3_B_wea          : t_IL_36_1b;
  signal IL_L6PHIC_neg2S_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_3_B_din         : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIC_neg2S_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHID_neg2S_3_B_start                   : std_logic;
  signal IL_L6PHID_neg2S_3_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHID_neg2S_3_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHID_neg2S_3_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHID_neg2S_3_B_wea          : t_IL_36_1b;
  signal IL_L6PHID_neg2S_3_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHID_neg2S_3_B_din         : t_IL_36_DATA;
  signal IL_L6PHID_neg2S_3_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHID_neg2S_3_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHID_neg2S_3_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHID_neg2S_3_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIA_neg2S_4_A_start                   : std_logic;
  signal IL_L6PHIA_neg2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIA_neg2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIA_neg2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIA_neg2S_4_A_wea          : t_IL_36_1b;
  signal IL_L6PHIA_neg2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIA_neg2S_4_A_din         : t_IL_36_DATA;
  signal IL_L6PHIA_neg2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIA_neg2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIA_neg2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIA_neg2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIB_neg2S_4_A_start                   : std_logic;
  signal IL_L6PHIB_neg2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIB_neg2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_4_A_wea          : t_IL_36_1b;
  signal IL_L6PHIB_neg2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_4_A_din         : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIB_neg2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIB_neg2S_4_B_start                   : std_logic;
  signal IL_L6PHIB_neg2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIB_neg2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_4_B_wea          : t_IL_36_1b;
  signal IL_L6PHIB_neg2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_4_B_din         : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIB_neg2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIB_neg2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIB_neg2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHIC_neg2S_4_B_start                   : std_logic;
  signal IL_L6PHIC_neg2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHIC_neg2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_4_B_wea          : t_IL_36_1b;
  signal IL_L6PHIC_neg2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_4_B_din         : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHIC_neg2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHIC_neg2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHIC_neg2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_L6PHID_neg2S_4_B_start                   : std_logic;
  signal IL_L6PHID_neg2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_L6PHID_neg2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_L6PHID_neg2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_L6PHID_neg2S_4_B_wea          : t_IL_36_1b;
  signal IL_L6PHID_neg2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_L6PHID_neg2S_4_B_din         : t_IL_36_DATA;
  signal IL_L6PHID_neg2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_L6PHID_neg2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_L6PHID_neg2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_L6PHID_neg2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIA_neg2S_4_A_start                   : std_logic;
  signal IL_D3PHIA_neg2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIA_neg2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIA_neg2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIA_neg2S_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIA_neg2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIA_neg2S_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIA_neg2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIA_neg2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIA_neg2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIA_neg2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_neg2S_4_A_start                   : std_logic;
  signal IL_D3PHIB_neg2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_neg2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_neg2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_neg2S_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIB_neg2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_neg2S_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIB_neg2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_neg2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_neg2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_neg2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIB_neg2S_4_B_start                   : std_logic;
  signal IL_D3PHIB_neg2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIB_neg2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIB_neg2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIB_neg2S_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIB_neg2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIB_neg2S_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIB_neg2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIB_neg2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIB_neg2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIB_neg2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_neg2S_4_A_start                   : std_logic;
  signal IL_D3PHIC_neg2S_4_A_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_neg2S_4_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_neg2S_4_A_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_neg2S_4_A_wea          : t_IL_36_1b;
  signal IL_D3PHIC_neg2S_4_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_neg2S_4_A_din         : t_IL_36_DATA;
  signal IL_D3PHIC_neg2S_4_A_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_neg2S_4_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_neg2S_4_A_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_neg2S_4_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHIC_neg2S_4_B_start                   : std_logic;
  signal IL_D3PHIC_neg2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHIC_neg2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHIC_neg2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHIC_neg2S_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHIC_neg2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHIC_neg2S_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHIC_neg2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHIC_neg2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHIC_neg2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHIC_neg2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D3PHID_neg2S_4_B_start                   : std_logic;
  signal IL_D3PHID_neg2S_4_B_wea_delay          : t_IL_36_1b;
  signal IL_D3PHID_neg2S_4_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D3PHID_neg2S_4_B_din_delay         : t_IL_36_DATA;
  signal IL_D3PHID_neg2S_4_B_wea          : t_IL_36_1b;
  signal IL_D3PHID_neg2S_4_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D3PHID_neg2S_4_B_din         : t_IL_36_DATA;
  signal IL_D3PHID_neg2S_4_B_enb          : t_IL_36_1b := '1';
  signal IL_D3PHID_neg2S_4_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D3PHID_neg2S_4_B_V_dout        : t_IL_36_DATA;
  signal IL_D3PHID_neg2S_4_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIA_neg2S_5_A_start                   : std_logic;
  signal IL_D1PHIA_neg2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIA_neg2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIA_neg2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIA_neg2S_5_A_wea          : t_IL_36_1b;
  signal IL_D1PHIA_neg2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIA_neg2S_5_A_din         : t_IL_36_DATA;
  signal IL_D1PHIA_neg2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIA_neg2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIA_neg2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIA_neg2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_neg2S_5_A_start                   : std_logic;
  signal IL_D1PHIB_neg2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_neg2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_neg2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_neg2S_5_A_wea          : t_IL_36_1b;
  signal IL_D1PHIB_neg2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_neg2S_5_A_din         : t_IL_36_DATA;
  signal IL_D1PHIB_neg2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_neg2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_neg2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_neg2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIB_neg2S_5_B_start                   : std_logic;
  signal IL_D1PHIB_neg2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIB_neg2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIB_neg2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIB_neg2S_5_B_wea          : t_IL_36_1b;
  signal IL_D1PHIB_neg2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIB_neg2S_5_B_din         : t_IL_36_DATA;
  signal IL_D1PHIB_neg2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIB_neg2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIB_neg2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIB_neg2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_neg2S_5_A_start                   : std_logic;
  signal IL_D1PHIC_neg2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_neg2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_neg2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_neg2S_5_A_wea          : t_IL_36_1b;
  signal IL_D1PHIC_neg2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_neg2S_5_A_din         : t_IL_36_DATA;
  signal IL_D1PHIC_neg2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_neg2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_neg2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_neg2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHIC_neg2S_5_B_start                   : std_logic;
  signal IL_D1PHIC_neg2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHIC_neg2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHIC_neg2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHIC_neg2S_5_B_wea          : t_IL_36_1b;
  signal IL_D1PHIC_neg2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHIC_neg2S_5_B_din         : t_IL_36_DATA;
  signal IL_D1PHIC_neg2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHIC_neg2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHIC_neg2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHIC_neg2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D1PHID_neg2S_5_B_start                   : std_logic;
  signal IL_D1PHID_neg2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D1PHID_neg2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D1PHID_neg2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D1PHID_neg2S_5_B_wea          : t_IL_36_1b;
  signal IL_D1PHID_neg2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D1PHID_neg2S_5_B_din         : t_IL_36_DATA;
  signal IL_D1PHID_neg2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D1PHID_neg2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D1PHID_neg2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D1PHID_neg2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIA_neg2S_5_A_start                   : std_logic;
  signal IL_D4PHIA_neg2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIA_neg2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIA_neg2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIA_neg2S_5_A_wea          : t_IL_36_1b;
  signal IL_D4PHIA_neg2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIA_neg2S_5_A_din         : t_IL_36_DATA;
  signal IL_D4PHIA_neg2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIA_neg2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIA_neg2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIA_neg2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_neg2S_5_A_start                   : std_logic;
  signal IL_D4PHIB_neg2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_neg2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_neg2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_neg2S_5_A_wea          : t_IL_36_1b;
  signal IL_D4PHIB_neg2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_neg2S_5_A_din         : t_IL_36_DATA;
  signal IL_D4PHIB_neg2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_neg2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_neg2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_neg2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIB_neg2S_5_B_start                   : std_logic;
  signal IL_D4PHIB_neg2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIB_neg2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIB_neg2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIB_neg2S_5_B_wea          : t_IL_36_1b;
  signal IL_D4PHIB_neg2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIB_neg2S_5_B_din         : t_IL_36_DATA;
  signal IL_D4PHIB_neg2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIB_neg2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIB_neg2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIB_neg2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_neg2S_5_A_start                   : std_logic;
  signal IL_D4PHIC_neg2S_5_A_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_neg2S_5_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_neg2S_5_A_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_neg2S_5_A_wea          : t_IL_36_1b;
  signal IL_D4PHIC_neg2S_5_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_neg2S_5_A_din         : t_IL_36_DATA;
  signal IL_D4PHIC_neg2S_5_A_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_neg2S_5_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_neg2S_5_A_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_neg2S_5_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHIC_neg2S_5_B_start                   : std_logic;
  signal IL_D4PHIC_neg2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHIC_neg2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHIC_neg2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHIC_neg2S_5_B_wea          : t_IL_36_1b;
  signal IL_D4PHIC_neg2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHIC_neg2S_5_B_din         : t_IL_36_DATA;
  signal IL_D4PHIC_neg2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHIC_neg2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHIC_neg2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHIC_neg2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D4PHID_neg2S_5_B_start                   : std_logic;
  signal IL_D4PHID_neg2S_5_B_wea_delay          : t_IL_36_1b;
  signal IL_D4PHID_neg2S_5_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D4PHID_neg2S_5_B_din_delay         : t_IL_36_DATA;
  signal IL_D4PHID_neg2S_5_B_wea          : t_IL_36_1b;
  signal IL_D4PHID_neg2S_5_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D4PHID_neg2S_5_B_din         : t_IL_36_DATA;
  signal IL_D4PHID_neg2S_5_B_enb          : t_IL_36_1b := '1';
  signal IL_D4PHID_neg2S_5_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D4PHID_neg2S_5_B_V_dout        : t_IL_36_DATA;
  signal IL_D4PHID_neg2S_5_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIA_neg2S_6_A_start                   : std_logic;
  signal IL_D2PHIA_neg2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIA_neg2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIA_neg2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIA_neg2S_6_A_wea          : t_IL_36_1b;
  signal IL_D2PHIA_neg2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIA_neg2S_6_A_din         : t_IL_36_DATA;
  signal IL_D2PHIA_neg2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIA_neg2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIA_neg2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIA_neg2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_neg2S_6_A_start                   : std_logic;
  signal IL_D2PHIB_neg2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_neg2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_neg2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_neg2S_6_A_wea          : t_IL_36_1b;
  signal IL_D2PHIB_neg2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_neg2S_6_A_din         : t_IL_36_DATA;
  signal IL_D2PHIB_neg2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_neg2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_neg2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_neg2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIB_neg2S_6_B_start                   : std_logic;
  signal IL_D2PHIB_neg2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIB_neg2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIB_neg2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIB_neg2S_6_B_wea          : t_IL_36_1b;
  signal IL_D2PHIB_neg2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIB_neg2S_6_B_din         : t_IL_36_DATA;
  signal IL_D2PHIB_neg2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIB_neg2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIB_neg2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIB_neg2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_neg2S_6_A_start                   : std_logic;
  signal IL_D2PHIC_neg2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_neg2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_neg2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_neg2S_6_A_wea          : t_IL_36_1b;
  signal IL_D2PHIC_neg2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_neg2S_6_A_din         : t_IL_36_DATA;
  signal IL_D2PHIC_neg2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_neg2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_neg2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_neg2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHIC_neg2S_6_B_start                   : std_logic;
  signal IL_D2PHIC_neg2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHIC_neg2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHIC_neg2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHIC_neg2S_6_B_wea          : t_IL_36_1b;
  signal IL_D2PHIC_neg2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHIC_neg2S_6_B_din         : t_IL_36_DATA;
  signal IL_D2PHIC_neg2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHIC_neg2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHIC_neg2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHIC_neg2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D2PHID_neg2S_6_B_start                   : std_logic;
  signal IL_D2PHID_neg2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D2PHID_neg2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D2PHID_neg2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D2PHID_neg2S_6_B_wea          : t_IL_36_1b;
  signal IL_D2PHID_neg2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D2PHID_neg2S_6_B_din         : t_IL_36_DATA;
  signal IL_D2PHID_neg2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D2PHID_neg2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D2PHID_neg2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D2PHID_neg2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIA_neg2S_6_A_start                   : std_logic;
  signal IL_D5PHIA_neg2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIA_neg2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIA_neg2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIA_neg2S_6_A_wea          : t_IL_36_1b;
  signal IL_D5PHIA_neg2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIA_neg2S_6_A_din         : t_IL_36_DATA;
  signal IL_D5PHIA_neg2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIA_neg2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIA_neg2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIA_neg2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_neg2S_6_A_start                   : std_logic;
  signal IL_D5PHIB_neg2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_neg2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_neg2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_neg2S_6_A_wea          : t_IL_36_1b;
  signal IL_D5PHIB_neg2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_neg2S_6_A_din         : t_IL_36_DATA;
  signal IL_D5PHIB_neg2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_neg2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_neg2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_neg2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIB_neg2S_6_B_start                   : std_logic;
  signal IL_D5PHIB_neg2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIB_neg2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIB_neg2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIB_neg2S_6_B_wea          : t_IL_36_1b;
  signal IL_D5PHIB_neg2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIB_neg2S_6_B_din         : t_IL_36_DATA;
  signal IL_D5PHIB_neg2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIB_neg2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIB_neg2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIB_neg2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_neg2S_6_A_start                   : std_logic;
  signal IL_D5PHIC_neg2S_6_A_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_neg2S_6_A_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_neg2S_6_A_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_neg2S_6_A_wea          : t_IL_36_1b;
  signal IL_D5PHIC_neg2S_6_A_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_neg2S_6_A_din         : t_IL_36_DATA;
  signal IL_D5PHIC_neg2S_6_A_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_neg2S_6_A_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_neg2S_6_A_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_neg2S_6_A_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHIC_neg2S_6_B_start                   : std_logic;
  signal IL_D5PHIC_neg2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHIC_neg2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHIC_neg2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHIC_neg2S_6_B_wea          : t_IL_36_1b;
  signal IL_D5PHIC_neg2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHIC_neg2S_6_B_din         : t_IL_36_DATA;
  signal IL_D5PHIC_neg2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHIC_neg2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHIC_neg2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHIC_neg2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal IL_D5PHID_neg2S_6_B_start                   : std_logic;
  signal IL_D5PHID_neg2S_6_B_wea_delay          : t_IL_36_1b;
  signal IL_D5PHID_neg2S_6_B_writeaddr_delay   : t_IL_36_ADDR;
  signal IL_D5PHID_neg2S_6_B_din_delay         : t_IL_36_DATA;
  signal IL_D5PHID_neg2S_6_B_wea          : t_IL_36_1b;
  signal IL_D5PHID_neg2S_6_B_writeaddr   : t_IL_36_ADDR;
  signal IL_D5PHID_neg2S_6_B_din         : t_IL_36_DATA;
  signal IL_D5PHID_neg2S_6_B_enb          : t_IL_36_1b := '1';
  signal IL_D5PHID_neg2S_6_B_V_readaddr    : t_IL_36_ADDR;
  signal IL_D5PHID_neg2S_6_B_V_dout        : t_IL_36_DATA;
  signal IL_D5PHID_neg2S_6_B_AV_dout_nent  : t_IL_36_NENT; -- (#page)
  signal AS_L1PHIAn1_start                   : std_logic;
  signal AS_L1PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIAn1_wea          : t_AS_36_1b;
  signal AS_L1PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIAn1_din         : t_AS_36_DATA;
  signal AS_L1PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIBn1_start                   : std_logic;
  signal AS_L1PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIBn1_wea          : t_AS_36_1b;
  signal AS_L1PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIBn1_din         : t_AS_36_DATA;
  signal AS_L1PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHICn1_start                   : std_logic;
  signal AS_L1PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHICn1_wea          : t_AS_36_1b;
  signal AS_L1PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHICn1_din         : t_AS_36_DATA;
  signal AS_L1PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIDn1_start                   : std_logic;
  signal AS_L1PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIDn1_wea          : t_AS_36_1b;
  signal AS_L1PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIDn1_din         : t_AS_36_DATA;
  signal AS_L1PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIEn1_start                   : std_logic;
  signal AS_L1PHIEn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIEn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIEn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIEn1_wea          : t_AS_36_1b;
  signal AS_L1PHIEn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIEn1_din         : t_AS_36_DATA;
  signal AS_L1PHIEn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHIEn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHIEn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHIEn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIFn1_start                   : std_logic;
  signal AS_L1PHIFn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIFn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIFn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIFn1_wea          : t_AS_36_1b;
  signal AS_L1PHIFn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIFn1_din         : t_AS_36_DATA;
  signal AS_L1PHIFn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHIFn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHIFn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHIFn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIGn1_start                   : std_logic;
  signal AS_L1PHIGn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIGn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIGn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIGn1_wea          : t_AS_36_1b;
  signal AS_L1PHIGn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIGn1_din         : t_AS_36_DATA;
  signal AS_L1PHIGn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHIGn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHIGn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHIGn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIHn1_start                   : std_logic;
  signal AS_L1PHIHn1_wea_delay          : t_AS_36_1b;
  signal AS_L1PHIHn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L1PHIHn1_din_delay         : t_AS_36_DATA;
  signal AS_L1PHIHn1_wea          : t_AS_36_1b;
  signal AS_L1PHIHn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L1PHIHn1_din         : t_AS_36_DATA;
  signal AS_L1PHIHn1_enb          : t_AS_36_1b := '1';
  --signal AS_L1PHIHn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L1PHIHn1_V_dout        : t_AS_36_DATA;
  --signal AS_L1PHIHn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIAn1_start                   : std_logic;
  signal AS_L2PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIAn1_wea          : t_AS_36_1b;
  signal AS_L2PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIAn1_din         : t_AS_36_DATA;
  signal AS_L2PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_L2PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L2PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_L2PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIBn1_start                   : std_logic;
  signal AS_L2PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIBn1_wea          : t_AS_36_1b;
  signal AS_L2PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIBn1_din         : t_AS_36_DATA;
  signal AS_L2PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_L2PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L2PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_L2PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHICn1_start                   : std_logic;
  signal AS_L2PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_L2PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_L2PHICn1_wea          : t_AS_36_1b;
  signal AS_L2PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHICn1_din         : t_AS_36_DATA;
  signal AS_L2PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_L2PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L2PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_L2PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIDn1_start                   : std_logic;
  signal AS_L2PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIDn1_wea          : t_AS_36_1b;
  signal AS_L2PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIDn1_din         : t_AS_36_DATA;
  signal AS_L2PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_L2PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L2PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_L2PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIAn1_start                   : std_logic;
  signal AS_L3PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIAn1_wea          : t_AS_36_1b;
  signal AS_L3PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIAn1_din         : t_AS_36_DATA;
  signal AS_L3PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_L3PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L3PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_L3PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIBn1_start                   : std_logic;
  signal AS_L3PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIBn1_wea          : t_AS_36_1b;
  signal AS_L3PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIBn1_din         : t_AS_36_DATA;
  signal AS_L3PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_L3PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L3PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_L3PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHICn1_start                   : std_logic;
  signal AS_L3PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_L3PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_L3PHICn1_wea          : t_AS_36_1b;
  signal AS_L3PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHICn1_din         : t_AS_36_DATA;
  signal AS_L3PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_L3PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L3PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_L3PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIDn1_start                   : std_logic;
  signal AS_L3PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIDn1_wea          : t_AS_36_1b;
  signal AS_L3PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIDn1_din         : t_AS_36_DATA;
  signal AS_L3PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_L3PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L3PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_L3PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIAn1_start                   : std_logic;
  signal AS_L4PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIAn1_wea          : t_AS_36_1b;
  signal AS_L4PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIAn1_din         : t_AS_36_DATA;
  signal AS_L4PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_L4PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L4PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_L4PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIBn1_start                   : std_logic;
  signal AS_L4PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIBn1_wea          : t_AS_36_1b;
  signal AS_L4PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIBn1_din         : t_AS_36_DATA;
  signal AS_L4PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_L4PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L4PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_L4PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHICn1_start                   : std_logic;
  signal AS_L4PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_L4PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_L4PHICn1_wea          : t_AS_36_1b;
  signal AS_L4PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHICn1_din         : t_AS_36_DATA;
  signal AS_L4PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_L4PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L4PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_L4PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIDn1_start                   : std_logic;
  signal AS_L4PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIDn1_wea          : t_AS_36_1b;
  signal AS_L4PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIDn1_din         : t_AS_36_DATA;
  signal AS_L4PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_L4PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L4PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_L4PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIAn1_start                   : std_logic;
  signal AS_L5PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIAn1_wea          : t_AS_36_1b;
  signal AS_L5PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHIAn1_din         : t_AS_36_DATA;
  signal AS_L5PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_L5PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L5PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_L5PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIBn1_start                   : std_logic;
  signal AS_L5PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIBn1_wea          : t_AS_36_1b;
  signal AS_L5PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHIBn1_din         : t_AS_36_DATA;
  signal AS_L5PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_L5PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L5PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_L5PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHICn1_start                   : std_logic;
  signal AS_L5PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_L5PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_L5PHICn1_wea          : t_AS_36_1b;
  signal AS_L5PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHICn1_din         : t_AS_36_DATA;
  signal AS_L5PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_L5PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L5PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_L5PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L5PHIDn1_start                   : std_logic;
  signal AS_L5PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_L5PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L5PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_L5PHIDn1_wea          : t_AS_36_1b;
  signal AS_L5PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L5PHIDn1_din         : t_AS_36_DATA;
  signal AS_L5PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_L5PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L5PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_L5PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIAn1_start                   : std_logic;
  signal AS_L6PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIAn1_wea          : t_AS_36_1b;
  signal AS_L6PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIAn1_din         : t_AS_36_DATA;
  signal AS_L6PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_L6PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L6PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_L6PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIBn1_start                   : std_logic;
  signal AS_L6PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIBn1_wea          : t_AS_36_1b;
  signal AS_L6PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIBn1_din         : t_AS_36_DATA;
  signal AS_L6PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_L6PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L6PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_L6PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHICn1_start                   : std_logic;
  signal AS_L6PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_L6PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_L6PHICn1_wea          : t_AS_36_1b;
  signal AS_L6PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHICn1_din         : t_AS_36_DATA;
  signal AS_L6PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_L6PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L6PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_L6PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIDn1_start                   : std_logic;
  signal AS_L6PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIDn1_wea          : t_AS_36_1b;
  signal AS_L6PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIDn1_din         : t_AS_36_DATA;
  signal AS_L6PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_L6PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_L6PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_L6PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIAn1_start                   : std_logic;
  signal AS_D1PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIAn1_wea          : t_AS_36_1b;
  signal AS_D1PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIAn1_din         : t_AS_36_DATA;
  signal AS_D1PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_D1PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D1PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_D1PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIBn1_start                   : std_logic;
  signal AS_D1PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIBn1_wea          : t_AS_36_1b;
  signal AS_D1PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIBn1_din         : t_AS_36_DATA;
  signal AS_D1PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_D1PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D1PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_D1PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHICn1_start                   : std_logic;
  signal AS_D1PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_D1PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_D1PHICn1_wea          : t_AS_36_1b;
  signal AS_D1PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHICn1_din         : t_AS_36_DATA;
  signal AS_D1PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_D1PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D1PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_D1PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIDn1_start                   : std_logic;
  signal AS_D1PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIDn1_wea          : t_AS_36_1b;
  signal AS_D1PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIDn1_din         : t_AS_36_DATA;
  signal AS_D1PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_D1PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D1PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_D1PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIAn1_start                   : std_logic;
  signal AS_D2PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIAn1_wea          : t_AS_36_1b;
  signal AS_D2PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIAn1_din         : t_AS_36_DATA;
  signal AS_D2PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_D2PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D2PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_D2PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIBn1_start                   : std_logic;
  signal AS_D2PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIBn1_wea          : t_AS_36_1b;
  signal AS_D2PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIBn1_din         : t_AS_36_DATA;
  signal AS_D2PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_D2PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D2PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_D2PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHICn1_start                   : std_logic;
  signal AS_D2PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_D2PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_D2PHICn1_wea          : t_AS_36_1b;
  signal AS_D2PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHICn1_din         : t_AS_36_DATA;
  signal AS_D2PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_D2PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D2PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_D2PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIDn1_start                   : std_logic;
  signal AS_D2PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIDn1_wea          : t_AS_36_1b;
  signal AS_D2PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIDn1_din         : t_AS_36_DATA;
  signal AS_D2PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_D2PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D2PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_D2PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIAn1_start                   : std_logic;
  signal AS_D3PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIAn1_wea          : t_AS_36_1b;
  signal AS_D3PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHIAn1_din         : t_AS_36_DATA;
  signal AS_D3PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_D3PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D3PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_D3PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIBn1_start                   : std_logic;
  signal AS_D3PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIBn1_wea          : t_AS_36_1b;
  signal AS_D3PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHIBn1_din         : t_AS_36_DATA;
  signal AS_D3PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_D3PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D3PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_D3PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHICn1_start                   : std_logic;
  signal AS_D3PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_D3PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_D3PHICn1_wea          : t_AS_36_1b;
  signal AS_D3PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHICn1_din         : t_AS_36_DATA;
  signal AS_D3PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_D3PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D3PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_D3PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D3PHIDn1_start                   : std_logic;
  signal AS_D3PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_D3PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D3PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_D3PHIDn1_wea          : t_AS_36_1b;
  signal AS_D3PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D3PHIDn1_din         : t_AS_36_DATA;
  signal AS_D3PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_D3PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D3PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_D3PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIAn1_start                   : std_logic;
  signal AS_D4PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIAn1_wea          : t_AS_36_1b;
  signal AS_D4PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIAn1_din         : t_AS_36_DATA;
  signal AS_D4PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_D4PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D4PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_D4PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIBn1_start                   : std_logic;
  signal AS_D4PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIBn1_wea          : t_AS_36_1b;
  signal AS_D4PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIBn1_din         : t_AS_36_DATA;
  signal AS_D4PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_D4PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D4PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_D4PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHICn1_start                   : std_logic;
  signal AS_D4PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_D4PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_D4PHICn1_wea          : t_AS_36_1b;
  signal AS_D4PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHICn1_din         : t_AS_36_DATA;
  signal AS_D4PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_D4PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D4PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_D4PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIDn1_start                   : std_logic;
  signal AS_D4PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIDn1_wea          : t_AS_36_1b;
  signal AS_D4PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIDn1_din         : t_AS_36_DATA;
  signal AS_D4PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_D4PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D4PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_D4PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIAn1_start                   : std_logic;
  signal AS_D5PHIAn1_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIAn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIAn1_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIAn1_wea          : t_AS_36_1b;
  signal AS_D5PHIAn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHIAn1_din         : t_AS_36_DATA;
  signal AS_D5PHIAn1_enb          : t_AS_36_1b := '1';
  --signal AS_D5PHIAn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D5PHIAn1_V_dout        : t_AS_36_DATA;
  --signal AS_D5PHIAn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIBn1_start                   : std_logic;
  signal AS_D5PHIBn1_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIBn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIBn1_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIBn1_wea          : t_AS_36_1b;
  signal AS_D5PHIBn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHIBn1_din         : t_AS_36_DATA;
  signal AS_D5PHIBn1_enb          : t_AS_36_1b := '1';
  --signal AS_D5PHIBn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D5PHIBn1_V_dout        : t_AS_36_DATA;
  --signal AS_D5PHIBn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHICn1_start                   : std_logic;
  signal AS_D5PHICn1_wea_delay          : t_AS_36_1b;
  signal AS_D5PHICn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHICn1_din_delay         : t_AS_36_DATA;
  signal AS_D5PHICn1_wea          : t_AS_36_1b;
  signal AS_D5PHICn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHICn1_din         : t_AS_36_DATA;
  signal AS_D5PHICn1_enb          : t_AS_36_1b := '1';
  --signal AS_D5PHICn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D5PHICn1_V_dout        : t_AS_36_DATA;
  --signal AS_D5PHICn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D5PHIDn1_start                   : std_logic;
  signal AS_D5PHIDn1_wea_delay          : t_AS_36_1b;
  signal AS_D5PHIDn1_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D5PHIDn1_din_delay         : t_AS_36_DATA;
  signal AS_D5PHIDn1_wea          : t_AS_36_1b;
  signal AS_D5PHIDn1_writeaddr   : t_AS_36_ADDR;
  signal AS_D5PHIDn1_din         : t_AS_36_DATA;
  signal AS_D5PHIDn1_enb          : t_AS_36_1b := '1';
  --signal AS_D5PHIDn1_V_readaddr    : t_AS_36_ADDR;
  --signal AS_D5PHIDn1_V_dout        : t_AS_36_DATA;
  --signal AS_D5PHIDn1_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIA_B_L1A_start                   : std_logic;
  signal AS_L2PHIA_B_L1A_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIA_B_L1A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1A_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1A_wea          : t_AS_36_1b;
  signal AS_L2PHIA_B_L1A_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1A_din         : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1A_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIA_B_L1A_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1A_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIA_B_L1B_start                   : std_logic;
  signal AS_L2PHIA_B_L1B_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIA_B_L1B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1B_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1B_wea          : t_AS_36_1b;
  signal AS_L2PHIA_B_L1B_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1B_din         : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1B_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIA_B_L1B_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1B_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIA_B_L1C_start                   : std_logic;
  signal AS_L2PHIA_B_L1C_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIA_B_L1C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1C_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1C_wea          : t_AS_36_1b;
  signal AS_L2PHIA_B_L1C_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1C_din         : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1C_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIA_B_L1C_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIA_B_L1C_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIA_B_L1C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIB_B_L1D_start                   : std_logic;
  signal AS_L2PHIB_B_L1D_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIB_B_L1D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1D_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1D_wea          : t_AS_36_1b;
  signal AS_L2PHIB_B_L1D_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1D_din         : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1D_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIB_B_L1D_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1D_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIB_B_L1E_start                   : std_logic;
  signal AS_L2PHIB_B_L1E_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIB_B_L1E_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1E_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1E_wea          : t_AS_36_1b;
  signal AS_L2PHIB_B_L1E_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1E_din         : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1E_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIB_B_L1E_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1E_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1E_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIB_B_L1F_start                   : std_logic;
  signal AS_L2PHIB_B_L1F_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIB_B_L1F_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1F_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1F_wea          : t_AS_36_1b;
  signal AS_L2PHIB_B_L1F_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1F_din         : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1F_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIB_B_L1F_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIB_B_L1F_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIB_B_L1F_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIC_B_L1G_start                   : std_logic;
  signal AS_L2PHIC_B_L1G_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIC_B_L1G_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1G_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1G_wea          : t_AS_36_1b;
  signal AS_L2PHIC_B_L1G_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1G_din         : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1G_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIC_B_L1G_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1G_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1G_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIC_B_L1H_start                   : std_logic;
  signal AS_L2PHIC_B_L1H_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIC_B_L1H_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1H_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1H_wea          : t_AS_36_1b;
  signal AS_L2PHIC_B_L1H_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1H_din         : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1H_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIC_B_L1H_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1H_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1H_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHIC_B_L1I_start                   : std_logic;
  signal AS_L2PHIC_B_L1I_wea_delay          : t_AS_36_1b;
  signal AS_L2PHIC_B_L1I_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1I_din_delay         : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1I_wea          : t_AS_36_1b;
  signal AS_L2PHIC_B_L1I_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1I_din         : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1I_enb          : t_AS_36_1b := '1';
  signal AS_L2PHIC_B_L1I_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHIC_B_L1I_V_dout        : t_AS_36_DATA;
  signal AS_L2PHIC_B_L1I_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHID_B_L1J_start                   : std_logic;
  signal AS_L2PHID_B_L1J_wea_delay          : t_AS_36_1b;
  signal AS_L2PHID_B_L1J_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1J_din_delay         : t_AS_36_DATA;
  signal AS_L2PHID_B_L1J_wea          : t_AS_36_1b;
  signal AS_L2PHID_B_L1J_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1J_din         : t_AS_36_DATA;
  signal AS_L2PHID_B_L1J_enb          : t_AS_36_1b := '1';
  signal AS_L2PHID_B_L1J_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1J_V_dout        : t_AS_36_DATA;
  signal AS_L2PHID_B_L1J_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHID_B_L1K_start                   : std_logic;
  signal AS_L2PHID_B_L1K_wea_delay          : t_AS_36_1b;
  signal AS_L2PHID_B_L1K_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1K_din_delay         : t_AS_36_DATA;
  signal AS_L2PHID_B_L1K_wea          : t_AS_36_1b;
  signal AS_L2PHID_B_L1K_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1K_din         : t_AS_36_DATA;
  signal AS_L2PHID_B_L1K_enb          : t_AS_36_1b := '1';
  signal AS_L2PHID_B_L1K_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1K_V_dout        : t_AS_36_DATA;
  signal AS_L2PHID_B_L1K_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L2PHID_B_L1L_start                   : std_logic;
  signal AS_L2PHID_B_L1L_wea_delay          : t_AS_36_1b;
  signal AS_L2PHID_B_L1L_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1L_din_delay         : t_AS_36_DATA;
  signal AS_L2PHID_B_L1L_wea          : t_AS_36_1b;
  signal AS_L2PHID_B_L1L_writeaddr   : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1L_din         : t_AS_36_DATA;
  signal AS_L2PHID_B_L1L_enb          : t_AS_36_1b := '1';
  signal AS_L2PHID_B_L1L_V_readaddr    : t_AS_36_ADDR;
  signal AS_L2PHID_B_L1L_V_dout        : t_AS_36_DATA;
  signal AS_L2PHID_B_L1L_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIA_B_L2A_start                   : std_logic;
  signal AS_L3PHIA_B_L2A_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIA_B_L2A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIA_B_L2A_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIA_B_L2A_wea          : t_AS_36_1b;
  signal AS_L3PHIA_B_L2A_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIA_B_L2A_din         : t_AS_36_DATA;
  signal AS_L3PHIA_B_L2A_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIA_B_L2A_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIA_B_L2A_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIA_B_L2A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIB_B_L2B_start                   : std_logic;
  signal AS_L3PHIB_B_L2B_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIB_B_L2B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIB_B_L2B_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIB_B_L2B_wea          : t_AS_36_1b;
  signal AS_L3PHIB_B_L2B_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIB_B_L2B_din         : t_AS_36_DATA;
  signal AS_L3PHIB_B_L2B_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIB_B_L2B_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIB_B_L2B_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIB_B_L2B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHIC_B_L2C_start                   : std_logic;
  signal AS_L3PHIC_B_L2C_wea_delay          : t_AS_36_1b;
  signal AS_L3PHIC_B_L2C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHIC_B_L2C_din_delay         : t_AS_36_DATA;
  signal AS_L3PHIC_B_L2C_wea          : t_AS_36_1b;
  signal AS_L3PHIC_B_L2C_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHIC_B_L2C_din         : t_AS_36_DATA;
  signal AS_L3PHIC_B_L2C_enb          : t_AS_36_1b := '1';
  signal AS_L3PHIC_B_L2C_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHIC_B_L2C_V_dout        : t_AS_36_DATA;
  signal AS_L3PHIC_B_L2C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L3PHID_B_L2D_start                   : std_logic;
  signal AS_L3PHID_B_L2D_wea_delay          : t_AS_36_1b;
  signal AS_L3PHID_B_L2D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L3PHID_B_L2D_din_delay         : t_AS_36_DATA;
  signal AS_L3PHID_B_L2D_wea          : t_AS_36_1b;
  signal AS_L3PHID_B_L2D_writeaddr   : t_AS_36_ADDR;
  signal AS_L3PHID_B_L2D_din         : t_AS_36_DATA;
  signal AS_L3PHID_B_L2D_enb          : t_AS_36_1b := '1';
  signal AS_L3PHID_B_L2D_V_readaddr    : t_AS_36_ADDR;
  signal AS_L3PHID_B_L2D_V_dout        : t_AS_36_DATA;
  signal AS_L3PHID_B_L2D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIA_B_L3A_start                   : std_logic;
  signal AS_L4PHIA_B_L3A_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIA_B_L3A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIA_B_L3A_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIA_B_L3A_wea          : t_AS_36_1b;
  signal AS_L4PHIA_B_L3A_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIA_B_L3A_din         : t_AS_36_DATA;
  signal AS_L4PHIA_B_L3A_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIA_B_L3A_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIA_B_L3A_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIA_B_L3A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIB_B_L3B_start                   : std_logic;
  signal AS_L4PHIB_B_L3B_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIB_B_L3B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIB_B_L3B_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIB_B_L3B_wea          : t_AS_36_1b;
  signal AS_L4PHIB_B_L3B_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIB_B_L3B_din         : t_AS_36_DATA;
  signal AS_L4PHIB_B_L3B_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIB_B_L3B_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIB_B_L3B_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIB_B_L3B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHIC_B_L3C_start                   : std_logic;
  signal AS_L4PHIC_B_L3C_wea_delay          : t_AS_36_1b;
  signal AS_L4PHIC_B_L3C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHIC_B_L3C_din_delay         : t_AS_36_DATA;
  signal AS_L4PHIC_B_L3C_wea          : t_AS_36_1b;
  signal AS_L4PHIC_B_L3C_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHIC_B_L3C_din         : t_AS_36_DATA;
  signal AS_L4PHIC_B_L3C_enb          : t_AS_36_1b := '1';
  signal AS_L4PHIC_B_L3C_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHIC_B_L3C_V_dout        : t_AS_36_DATA;
  signal AS_L4PHIC_B_L3C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L4PHID_B_L3D_start                   : std_logic;
  signal AS_L4PHID_B_L3D_wea_delay          : t_AS_36_1b;
  signal AS_L4PHID_B_L3D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L4PHID_B_L3D_din_delay         : t_AS_36_DATA;
  signal AS_L4PHID_B_L3D_wea          : t_AS_36_1b;
  signal AS_L4PHID_B_L3D_writeaddr   : t_AS_36_ADDR;
  signal AS_L4PHID_B_L3D_din         : t_AS_36_DATA;
  signal AS_L4PHID_B_L3D_enb          : t_AS_36_1b := '1';
  signal AS_L4PHID_B_L3D_V_readaddr    : t_AS_36_ADDR;
  signal AS_L4PHID_B_L3D_V_dout        : t_AS_36_DATA;
  signal AS_L4PHID_B_L3D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIA_B_L5A_start                   : std_logic;
  signal AS_L6PHIA_B_L5A_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIA_B_L5A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIA_B_L5A_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIA_B_L5A_wea          : t_AS_36_1b;
  signal AS_L6PHIA_B_L5A_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIA_B_L5A_din         : t_AS_36_DATA;
  signal AS_L6PHIA_B_L5A_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIA_B_L5A_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIA_B_L5A_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIA_B_L5A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIB_B_L5B_start                   : std_logic;
  signal AS_L6PHIB_B_L5B_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIB_B_L5B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIB_B_L5B_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIB_B_L5B_wea          : t_AS_36_1b;
  signal AS_L6PHIB_B_L5B_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIB_B_L5B_din         : t_AS_36_DATA;
  signal AS_L6PHIB_B_L5B_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIB_B_L5B_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIB_B_L5B_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIB_B_L5B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHIC_B_L5C_start                   : std_logic;
  signal AS_L6PHIC_B_L5C_wea_delay          : t_AS_36_1b;
  signal AS_L6PHIC_B_L5C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHIC_B_L5C_din_delay         : t_AS_36_DATA;
  signal AS_L6PHIC_B_L5C_wea          : t_AS_36_1b;
  signal AS_L6PHIC_B_L5C_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHIC_B_L5C_din         : t_AS_36_DATA;
  signal AS_L6PHIC_B_L5C_enb          : t_AS_36_1b := '1';
  signal AS_L6PHIC_B_L5C_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHIC_B_L5C_V_dout        : t_AS_36_DATA;
  signal AS_L6PHIC_B_L5C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L6PHID_B_L5D_start                   : std_logic;
  signal AS_L6PHID_B_L5D_wea_delay          : t_AS_36_1b;
  signal AS_L6PHID_B_L5D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_L6PHID_B_L5D_din_delay         : t_AS_36_DATA;
  signal AS_L6PHID_B_L5D_wea          : t_AS_36_1b;
  signal AS_L6PHID_B_L5D_writeaddr   : t_AS_36_ADDR;
  signal AS_L6PHID_B_L5D_din         : t_AS_36_DATA;
  signal AS_L6PHID_B_L5D_enb          : t_AS_36_1b := '1';
  signal AS_L6PHID_B_L5D_V_readaddr    : t_AS_36_ADDR;
  signal AS_L6PHID_B_L5D_V_dout        : t_AS_36_DATA;
  signal AS_L6PHID_B_L5D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIA_O_L1A_start                   : std_logic;
  signal AS_D1PHIA_O_L1A_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIA_O_L1A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L1A_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIA_O_L1A_wea          : t_AS_36_1b;
  signal AS_D1PHIA_O_L1A_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L1A_din         : t_AS_36_DATA;
  signal AS_D1PHIA_O_L1A_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIA_O_L1A_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L1A_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIA_O_L1A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIA_O_L1B_start                   : std_logic;
  signal AS_D1PHIA_O_L1B_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIA_O_L1B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L1B_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIA_O_L1B_wea          : t_AS_36_1b;
  signal AS_D1PHIA_O_L1B_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L1B_din         : t_AS_36_DATA;
  signal AS_D1PHIA_O_L1B_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIA_O_L1B_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L1B_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIA_O_L1B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIA_O_L2A_start                   : std_logic;
  signal AS_D1PHIA_O_L2A_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIA_O_L2A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L2A_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIA_O_L2A_wea          : t_AS_36_1b;
  signal AS_D1PHIA_O_L2A_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L2A_din         : t_AS_36_DATA;
  signal AS_D1PHIA_O_L2A_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIA_O_L2A_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIA_O_L2A_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIA_O_L2A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIB_O_L1C_start                   : std_logic;
  signal AS_D1PHIB_O_L1C_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIB_O_L1C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L1C_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIB_O_L1C_wea          : t_AS_36_1b;
  signal AS_D1PHIB_O_L1C_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L1C_din         : t_AS_36_DATA;
  signal AS_D1PHIB_O_L1C_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIB_O_L1C_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L1C_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIB_O_L1C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIB_O_L1D_start                   : std_logic;
  signal AS_D1PHIB_O_L1D_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIB_O_L1D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L1D_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIB_O_L1D_wea          : t_AS_36_1b;
  signal AS_D1PHIB_O_L1D_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L1D_din         : t_AS_36_DATA;
  signal AS_D1PHIB_O_L1D_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIB_O_L1D_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L1D_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIB_O_L1D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIB_O_L2B_start                   : std_logic;
  signal AS_D1PHIB_O_L2B_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIB_O_L2B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L2B_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIB_O_L2B_wea          : t_AS_36_1b;
  signal AS_D1PHIB_O_L2B_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L2B_din         : t_AS_36_DATA;
  signal AS_D1PHIB_O_L2B_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIB_O_L2B_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIB_O_L2B_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIB_O_L2B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIC_O_L1E_start                   : std_logic;
  signal AS_D1PHIC_O_L1E_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIC_O_L1E_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L1E_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIC_O_L1E_wea          : t_AS_36_1b;
  signal AS_D1PHIC_O_L1E_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L1E_din         : t_AS_36_DATA;
  signal AS_D1PHIC_O_L1E_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIC_O_L1E_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L1E_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIC_O_L1E_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIC_O_L1F_start                   : std_logic;
  signal AS_D1PHIC_O_L1F_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIC_O_L1F_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L1F_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIC_O_L1F_wea          : t_AS_36_1b;
  signal AS_D1PHIC_O_L1F_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L1F_din         : t_AS_36_DATA;
  signal AS_D1PHIC_O_L1F_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIC_O_L1F_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L1F_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIC_O_L1F_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHIC_O_L2C_start                   : std_logic;
  signal AS_D1PHIC_O_L2C_wea_delay          : t_AS_36_1b;
  signal AS_D1PHIC_O_L2C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L2C_din_delay         : t_AS_36_DATA;
  signal AS_D1PHIC_O_L2C_wea          : t_AS_36_1b;
  signal AS_D1PHIC_O_L2C_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L2C_din         : t_AS_36_DATA;
  signal AS_D1PHIC_O_L2C_enb          : t_AS_36_1b := '1';
  signal AS_D1PHIC_O_L2C_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHIC_O_L2C_V_dout        : t_AS_36_DATA;
  signal AS_D1PHIC_O_L2C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHID_O_L1G_start                   : std_logic;
  signal AS_D1PHID_O_L1G_wea_delay          : t_AS_36_1b;
  signal AS_D1PHID_O_L1G_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHID_O_L1G_din_delay         : t_AS_36_DATA;
  signal AS_D1PHID_O_L1G_wea          : t_AS_36_1b;
  signal AS_D1PHID_O_L1G_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHID_O_L1G_din         : t_AS_36_DATA;
  signal AS_D1PHID_O_L1G_enb          : t_AS_36_1b := '1';
  signal AS_D1PHID_O_L1G_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHID_O_L1G_V_dout        : t_AS_36_DATA;
  signal AS_D1PHID_O_L1G_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHID_O_L1H_start                   : std_logic;
  signal AS_D1PHID_O_L1H_wea_delay          : t_AS_36_1b;
  signal AS_D1PHID_O_L1H_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHID_O_L1H_din_delay         : t_AS_36_DATA;
  signal AS_D1PHID_O_L1H_wea          : t_AS_36_1b;
  signal AS_D1PHID_O_L1H_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHID_O_L1H_din         : t_AS_36_DATA;
  signal AS_D1PHID_O_L1H_enb          : t_AS_36_1b := '1';
  signal AS_D1PHID_O_L1H_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHID_O_L1H_V_dout        : t_AS_36_DATA;
  signal AS_D1PHID_O_L1H_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D1PHID_O_L2D_start                   : std_logic;
  signal AS_D1PHID_O_L2D_wea_delay          : t_AS_36_1b;
  signal AS_D1PHID_O_L2D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D1PHID_O_L2D_din_delay         : t_AS_36_DATA;
  signal AS_D1PHID_O_L2D_wea          : t_AS_36_1b;
  signal AS_D1PHID_O_L2D_writeaddr   : t_AS_36_ADDR;
  signal AS_D1PHID_O_L2D_din         : t_AS_36_DATA;
  signal AS_D1PHID_O_L2D_enb          : t_AS_36_1b := '1';
  signal AS_D1PHID_O_L2D_V_readaddr    : t_AS_36_ADDR;
  signal AS_D1PHID_O_L2D_V_dout        : t_AS_36_DATA;
  signal AS_D1PHID_O_L2D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIA_D_D1A_start                   : std_logic;
  signal AS_D2PHIA_D_D1A_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIA_D_D1A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIA_D_D1A_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIA_D_D1A_wea          : t_AS_36_1b;
  signal AS_D2PHIA_D_D1A_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIA_D_D1A_din         : t_AS_36_DATA;
  signal AS_D2PHIA_D_D1A_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIA_D_D1A_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIA_D_D1A_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIA_D_D1A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIB_D_D1B_start                   : std_logic;
  signal AS_D2PHIB_D_D1B_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIB_D_D1B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIB_D_D1B_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIB_D_D1B_wea          : t_AS_36_1b;
  signal AS_D2PHIB_D_D1B_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIB_D_D1B_din         : t_AS_36_DATA;
  signal AS_D2PHIB_D_D1B_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIB_D_D1B_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIB_D_D1B_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIB_D_D1B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHIC_D_D1C_start                   : std_logic;
  signal AS_D2PHIC_D_D1C_wea_delay          : t_AS_36_1b;
  signal AS_D2PHIC_D_D1C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHIC_D_D1C_din_delay         : t_AS_36_DATA;
  signal AS_D2PHIC_D_D1C_wea          : t_AS_36_1b;
  signal AS_D2PHIC_D_D1C_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHIC_D_D1C_din         : t_AS_36_DATA;
  signal AS_D2PHIC_D_D1C_enb          : t_AS_36_1b := '1';
  signal AS_D2PHIC_D_D1C_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHIC_D_D1C_V_dout        : t_AS_36_DATA;
  signal AS_D2PHIC_D_D1C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D2PHID_D_D1D_start                   : std_logic;
  signal AS_D2PHID_D_D1D_wea_delay          : t_AS_36_1b;
  signal AS_D2PHID_D_D1D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D2PHID_D_D1D_din_delay         : t_AS_36_DATA;
  signal AS_D2PHID_D_D1D_wea          : t_AS_36_1b;
  signal AS_D2PHID_D_D1D_writeaddr   : t_AS_36_ADDR;
  signal AS_D2PHID_D_D1D_din         : t_AS_36_DATA;
  signal AS_D2PHID_D_D1D_enb          : t_AS_36_1b := '1';
  signal AS_D2PHID_D_D1D_V_readaddr    : t_AS_36_ADDR;
  signal AS_D2PHID_D_D1D_V_dout        : t_AS_36_DATA;
  signal AS_D2PHID_D_D1D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIA_D_D3A_start                   : std_logic;
  signal AS_D4PHIA_D_D3A_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIA_D_D3A_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIA_D_D3A_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIA_D_D3A_wea          : t_AS_36_1b;
  signal AS_D4PHIA_D_D3A_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIA_D_D3A_din         : t_AS_36_DATA;
  signal AS_D4PHIA_D_D3A_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIA_D_D3A_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIA_D_D3A_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIA_D_D3A_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIB_D_D3B_start                   : std_logic;
  signal AS_D4PHIB_D_D3B_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIB_D_D3B_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIB_D_D3B_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIB_D_D3B_wea          : t_AS_36_1b;
  signal AS_D4PHIB_D_D3B_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIB_D_D3B_din         : t_AS_36_DATA;
  signal AS_D4PHIB_D_D3B_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIB_D_D3B_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIB_D_D3B_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIB_D_D3B_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHIC_D_D3C_start                   : std_logic;
  signal AS_D4PHIC_D_D3C_wea_delay          : t_AS_36_1b;
  signal AS_D4PHIC_D_D3C_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHIC_D_D3C_din_delay         : t_AS_36_DATA;
  signal AS_D4PHIC_D_D3C_wea          : t_AS_36_1b;
  signal AS_D4PHIC_D_D3C_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHIC_D_D3C_din         : t_AS_36_DATA;
  signal AS_D4PHIC_D_D3C_enb          : t_AS_36_1b := '1';
  signal AS_D4PHIC_D_D3C_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHIC_D_D3C_V_dout        : t_AS_36_DATA;
  signal AS_D4PHIC_D_D3C_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_D4PHID_D_D3D_start                   : std_logic;
  signal AS_D4PHID_D_D3D_wea_delay          : t_AS_36_1b;
  signal AS_D4PHID_D_D3D_writeaddr_delay   : t_AS_36_ADDR;
  signal AS_D4PHID_D_D3D_din_delay         : t_AS_36_DATA;
  signal AS_D4PHID_D_D3D_wea          : t_AS_36_1b;
  signal AS_D4PHID_D_D3D_writeaddr   : t_AS_36_ADDR;
  signal AS_D4PHID_D_D3D_din         : t_AS_36_DATA;
  signal AS_D4PHID_D_D3D_enb          : t_AS_36_1b := '1';
  signal AS_D4PHID_D_D3D_V_readaddr    : t_AS_36_ADDR;
  signal AS_D4PHID_D_D3D_V_dout        : t_AS_36_DATA;
  signal AS_D4PHID_D_D3D_AV_dout_nent  : t_AS_36_NENT; -- (#page)
  signal AS_L1PHIA_BF_start                   : std_logic;
  signal AS_L1PHIA_BF_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIA_BF_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIA_BF_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIA_BF_wea          : t_AS_51_1b;
  signal AS_L1PHIA_BF_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIA_BF_din         : t_AS_51_DATA;
  signal AS_L1PHIA_BF_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIA_BF_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIA_BF_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIA_BF_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIA_BE_start                   : std_logic;
  signal AS_L1PHIA_BE_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIA_BE_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIA_BE_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIA_BE_wea          : t_AS_51_1b;
  signal AS_L1PHIA_BE_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIA_BE_din         : t_AS_51_DATA;
  signal AS_L1PHIA_BE_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIA_BE_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIA_BE_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIA_BE_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIA_OM_start                   : std_logic;
  signal AS_L1PHIA_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIA_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIA_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIA_OM_wea          : t_AS_51_1b;
  signal AS_L1PHIA_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIA_OM_din         : t_AS_51_DATA;
  signal AS_L1PHIA_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIA_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIA_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIA_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIB_BD_start                   : std_logic;
  signal AS_L1PHIB_BD_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIB_BD_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIB_BD_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIB_BD_wea          : t_AS_51_1b;
  signal AS_L1PHIB_BD_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIB_BD_din         : t_AS_51_DATA;
  signal AS_L1PHIB_BD_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIB_BD_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIB_BD_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIB_BD_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIB_BC_start                   : std_logic;
  signal AS_L1PHIB_BC_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIB_BC_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIB_BC_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIB_BC_wea          : t_AS_51_1b;
  signal AS_L1PHIB_BC_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIB_BC_din         : t_AS_51_DATA;
  signal AS_L1PHIB_BC_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIB_BC_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIB_BC_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIB_BC_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIB_BA_start                   : std_logic;
  signal AS_L1PHIB_BA_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIB_BA_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIB_BA_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIB_BA_wea          : t_AS_51_1b;
  signal AS_L1PHIB_BA_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIB_BA_din         : t_AS_51_DATA;
  signal AS_L1PHIB_BA_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIB_BA_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIB_BA_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIB_BA_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIB_OM_start                   : std_logic;
  signal AS_L1PHIB_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIB_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIB_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIB_OM_wea          : t_AS_51_1b;
  signal AS_L1PHIB_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIB_OM_din         : t_AS_51_DATA;
  signal AS_L1PHIB_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIB_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIB_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIB_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIB_OR_start                   : std_logic;
  signal AS_L1PHIB_OR_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIB_OR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIB_OR_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIB_OR_wea          : t_AS_51_1b;
  signal AS_L1PHIB_OR_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIB_OR_din         : t_AS_51_DATA;
  signal AS_L1PHIB_OR_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIB_OR_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIB_OR_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIB_OR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIC_BB_start                   : std_logic;
  signal AS_L1PHIC_BB_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIC_BB_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIC_BB_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIC_BB_wea          : t_AS_51_1b;
  signal AS_L1PHIC_BB_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIC_BB_din         : t_AS_51_DATA;
  signal AS_L1PHIC_BB_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIC_BB_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIC_BB_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIC_BB_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIC_BF_start                   : std_logic;
  signal AS_L1PHIC_BF_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIC_BF_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIC_BF_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIC_BF_wea          : t_AS_51_1b;
  signal AS_L1PHIC_BF_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIC_BF_din         : t_AS_51_DATA;
  signal AS_L1PHIC_BF_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIC_BF_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIC_BF_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIC_BF_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIC_BE_start                   : std_logic;
  signal AS_L1PHIC_BE_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIC_BE_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIC_BE_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIC_BE_wea          : t_AS_51_1b;
  signal AS_L1PHIC_BE_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIC_BE_din         : t_AS_51_DATA;
  signal AS_L1PHIC_BE_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIC_BE_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIC_BE_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIC_BE_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIC_OL_start                   : std_logic;
  signal AS_L1PHIC_OL_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIC_OL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIC_OL_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIC_OL_wea          : t_AS_51_1b;
  signal AS_L1PHIC_OL_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIC_OL_din         : t_AS_51_DATA;
  signal AS_L1PHIC_OL_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIC_OL_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIC_OL_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIC_OL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIC_OM_start                   : std_logic;
  signal AS_L1PHIC_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIC_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIC_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIC_OM_wea          : t_AS_51_1b;
  signal AS_L1PHIC_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIC_OM_din         : t_AS_51_DATA;
  signal AS_L1PHIC_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIC_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIC_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIC_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHID_BD_start                   : std_logic;
  signal AS_L1PHID_BD_wea_delay          : t_AS_51_1b;
  signal AS_L1PHID_BD_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHID_BD_din_delay         : t_AS_51_DATA;
  signal AS_L1PHID_BD_wea          : t_AS_51_1b;
  signal AS_L1PHID_BD_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHID_BD_din         : t_AS_51_DATA;
  signal AS_L1PHID_BD_enb          : t_AS_51_1b := '1';
  signal AS_L1PHID_BD_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHID_BD_V_dout        : t_AS_51_DATA;
  signal AS_L1PHID_BD_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHID_BC_start                   : std_logic;
  signal AS_L1PHID_BC_wea_delay          : t_AS_51_1b;
  signal AS_L1PHID_BC_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHID_BC_din_delay         : t_AS_51_DATA;
  signal AS_L1PHID_BC_wea          : t_AS_51_1b;
  signal AS_L1PHID_BC_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHID_BC_din         : t_AS_51_DATA;
  signal AS_L1PHID_BC_enb          : t_AS_51_1b := '1';
  signal AS_L1PHID_BC_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHID_BC_V_dout        : t_AS_51_DATA;
  signal AS_L1PHID_BC_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHID_BA_start                   : std_logic;
  signal AS_L1PHID_BA_wea_delay          : t_AS_51_1b;
  signal AS_L1PHID_BA_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHID_BA_din_delay         : t_AS_51_DATA;
  signal AS_L1PHID_BA_wea          : t_AS_51_1b;
  signal AS_L1PHID_BA_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHID_BA_din         : t_AS_51_DATA;
  signal AS_L1PHID_BA_enb          : t_AS_51_1b := '1';
  signal AS_L1PHID_BA_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHID_BA_V_dout        : t_AS_51_DATA;
  signal AS_L1PHID_BA_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHID_OM_start                   : std_logic;
  signal AS_L1PHID_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHID_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHID_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHID_OM_wea          : t_AS_51_1b;
  signal AS_L1PHID_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHID_OM_din         : t_AS_51_DATA;
  signal AS_L1PHID_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHID_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHID_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHID_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHID_OR_start                   : std_logic;
  signal AS_L1PHID_OR_wea_delay          : t_AS_51_1b;
  signal AS_L1PHID_OR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHID_OR_din_delay         : t_AS_51_DATA;
  signal AS_L1PHID_OR_wea          : t_AS_51_1b;
  signal AS_L1PHID_OR_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHID_OR_din         : t_AS_51_DATA;
  signal AS_L1PHID_OR_enb          : t_AS_51_1b := '1';
  signal AS_L1PHID_OR_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHID_OR_V_dout        : t_AS_51_DATA;
  signal AS_L1PHID_OR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIE_BB_start                   : std_logic;
  signal AS_L1PHIE_BB_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIE_BB_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIE_BB_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIE_BB_wea          : t_AS_51_1b;
  signal AS_L1PHIE_BB_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIE_BB_din         : t_AS_51_DATA;
  signal AS_L1PHIE_BB_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIE_BB_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIE_BB_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIE_BB_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIE_BF_start                   : std_logic;
  signal AS_L1PHIE_BF_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIE_BF_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIE_BF_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIE_BF_wea          : t_AS_51_1b;
  signal AS_L1PHIE_BF_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIE_BF_din         : t_AS_51_DATA;
  signal AS_L1PHIE_BF_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIE_BF_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIE_BF_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIE_BF_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIE_BE_start                   : std_logic;
  signal AS_L1PHIE_BE_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIE_BE_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIE_BE_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIE_BE_wea          : t_AS_51_1b;
  signal AS_L1PHIE_BE_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIE_BE_din         : t_AS_51_DATA;
  signal AS_L1PHIE_BE_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIE_BE_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIE_BE_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIE_BE_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIE_OL_start                   : std_logic;
  signal AS_L1PHIE_OL_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIE_OL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIE_OL_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIE_OL_wea          : t_AS_51_1b;
  signal AS_L1PHIE_OL_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIE_OL_din         : t_AS_51_DATA;
  signal AS_L1PHIE_OL_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIE_OL_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIE_OL_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIE_OL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIE_OM_start                   : std_logic;
  signal AS_L1PHIE_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIE_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIE_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIE_OM_wea          : t_AS_51_1b;
  signal AS_L1PHIE_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIE_OM_din         : t_AS_51_DATA;
  signal AS_L1PHIE_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIE_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIE_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIE_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIF_BD_start                   : std_logic;
  signal AS_L1PHIF_BD_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIF_BD_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIF_BD_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIF_BD_wea          : t_AS_51_1b;
  signal AS_L1PHIF_BD_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIF_BD_din         : t_AS_51_DATA;
  signal AS_L1PHIF_BD_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIF_BD_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIF_BD_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIF_BD_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIF_BC_start                   : std_logic;
  signal AS_L1PHIF_BC_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIF_BC_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIF_BC_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIF_BC_wea          : t_AS_51_1b;
  signal AS_L1PHIF_BC_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIF_BC_din         : t_AS_51_DATA;
  signal AS_L1PHIF_BC_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIF_BC_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIF_BC_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIF_BC_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIF_BA_start                   : std_logic;
  signal AS_L1PHIF_BA_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIF_BA_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIF_BA_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIF_BA_wea          : t_AS_51_1b;
  signal AS_L1PHIF_BA_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIF_BA_din         : t_AS_51_DATA;
  signal AS_L1PHIF_BA_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIF_BA_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIF_BA_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIF_BA_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIF_OM_start                   : std_logic;
  signal AS_L1PHIF_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIF_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIF_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIF_OM_wea          : t_AS_51_1b;
  signal AS_L1PHIF_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIF_OM_din         : t_AS_51_DATA;
  signal AS_L1PHIF_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIF_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIF_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIF_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIF_OR_start                   : std_logic;
  signal AS_L1PHIF_OR_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIF_OR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIF_OR_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIF_OR_wea          : t_AS_51_1b;
  signal AS_L1PHIF_OR_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIF_OR_din         : t_AS_51_DATA;
  signal AS_L1PHIF_OR_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIF_OR_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIF_OR_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIF_OR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIG_BB_start                   : std_logic;
  signal AS_L1PHIG_BB_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIG_BB_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIG_BB_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIG_BB_wea          : t_AS_51_1b;
  signal AS_L1PHIG_BB_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIG_BB_din         : t_AS_51_DATA;
  signal AS_L1PHIG_BB_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIG_BB_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIG_BB_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIG_BB_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIG_BF_start                   : std_logic;
  signal AS_L1PHIG_BF_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIG_BF_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIG_BF_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIG_BF_wea          : t_AS_51_1b;
  signal AS_L1PHIG_BF_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIG_BF_din         : t_AS_51_DATA;
  signal AS_L1PHIG_BF_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIG_BF_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIG_BF_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIG_BF_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIG_BE_start                   : std_logic;
  signal AS_L1PHIG_BE_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIG_BE_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIG_BE_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIG_BE_wea          : t_AS_51_1b;
  signal AS_L1PHIG_BE_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIG_BE_din         : t_AS_51_DATA;
  signal AS_L1PHIG_BE_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIG_BE_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIG_BE_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIG_BE_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIG_OL_start                   : std_logic;
  signal AS_L1PHIG_OL_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIG_OL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIG_OL_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIG_OL_wea          : t_AS_51_1b;
  signal AS_L1PHIG_OL_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIG_OL_din         : t_AS_51_DATA;
  signal AS_L1PHIG_OL_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIG_OL_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIG_OL_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIG_OL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIG_OM_start                   : std_logic;
  signal AS_L1PHIG_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIG_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIG_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIG_OM_wea          : t_AS_51_1b;
  signal AS_L1PHIG_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIG_OM_din         : t_AS_51_DATA;
  signal AS_L1PHIG_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIG_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIG_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIG_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIH_BD_start                   : std_logic;
  signal AS_L1PHIH_BD_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIH_BD_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIH_BD_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIH_BD_wea          : t_AS_51_1b;
  signal AS_L1PHIH_BD_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIH_BD_din         : t_AS_51_DATA;
  signal AS_L1PHIH_BD_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIH_BD_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIH_BD_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIH_BD_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIH_BC_start                   : std_logic;
  signal AS_L1PHIH_BC_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIH_BC_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIH_BC_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIH_BC_wea          : t_AS_51_1b;
  signal AS_L1PHIH_BC_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIH_BC_din         : t_AS_51_DATA;
  signal AS_L1PHIH_BC_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIH_BC_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIH_BC_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIH_BC_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L1PHIH_OM_start                   : std_logic;
  signal AS_L1PHIH_OM_wea_delay          : t_AS_51_1b;
  signal AS_L1PHIH_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L1PHIH_OM_din_delay         : t_AS_51_DATA;
  signal AS_L1PHIH_OM_wea          : t_AS_51_1b;
  signal AS_L1PHIH_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L1PHIH_OM_din         : t_AS_51_DATA;
  signal AS_L1PHIH_OM_enb          : t_AS_51_1b := '1';
  signal AS_L1PHIH_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L1PHIH_OM_V_dout        : t_AS_51_DATA;
  signal AS_L1PHIH_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIA_BM_start                   : std_logic;
  signal AS_L2PHIA_BM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIA_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIA_BM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIA_BM_wea          : t_AS_51_1b;
  signal AS_L2PHIA_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIA_BM_din         : t_AS_51_DATA;
  signal AS_L2PHIA_BM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIA_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIA_BM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIA_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIA_OM_start                   : std_logic;
  signal AS_L2PHIA_OM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIA_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIA_OM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIA_OM_wea          : t_AS_51_1b;
  signal AS_L2PHIA_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIA_OM_din         : t_AS_51_DATA;
  signal AS_L2PHIA_OM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIA_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIA_OM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIA_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIB_BM_start                   : std_logic;
  signal AS_L2PHIB_BM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIB_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIB_BM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIB_BM_wea          : t_AS_51_1b;
  signal AS_L2PHIB_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIB_BM_din         : t_AS_51_DATA;
  signal AS_L2PHIB_BM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIB_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIB_BM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIB_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIB_BR_start                   : std_logic;
  signal AS_L2PHIB_BR_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIB_BR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIB_BR_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIB_BR_wea          : t_AS_51_1b;
  signal AS_L2PHIB_BR_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIB_BR_din         : t_AS_51_DATA;
  signal AS_L2PHIB_BR_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIB_BR_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIB_BR_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIB_BR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIB_OM_start                   : std_logic;
  signal AS_L2PHIB_OM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIB_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIB_OM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIB_OM_wea          : t_AS_51_1b;
  signal AS_L2PHIB_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIB_OM_din         : t_AS_51_DATA;
  signal AS_L2PHIB_OM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIB_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIB_OM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIB_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIB_OR_start                   : std_logic;
  signal AS_L2PHIB_OR_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIB_OR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIB_OR_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIB_OR_wea          : t_AS_51_1b;
  signal AS_L2PHIB_OR_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIB_OR_din         : t_AS_51_DATA;
  signal AS_L2PHIB_OR_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIB_OR_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIB_OR_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIB_OR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIC_BL_start                   : std_logic;
  signal AS_L2PHIC_BL_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIC_BL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIC_BL_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIC_BL_wea          : t_AS_51_1b;
  signal AS_L2PHIC_BL_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIC_BL_din         : t_AS_51_DATA;
  signal AS_L2PHIC_BL_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIC_BL_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIC_BL_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIC_BL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIC_BM_start                   : std_logic;
  signal AS_L2PHIC_BM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIC_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIC_BM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIC_BM_wea          : t_AS_51_1b;
  signal AS_L2PHIC_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIC_BM_din         : t_AS_51_DATA;
  signal AS_L2PHIC_BM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIC_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIC_BM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIC_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIC_OL_start                   : std_logic;
  signal AS_L2PHIC_OL_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIC_OL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIC_OL_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIC_OL_wea          : t_AS_51_1b;
  signal AS_L2PHIC_OL_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIC_OL_din         : t_AS_51_DATA;
  signal AS_L2PHIC_OL_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIC_OL_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIC_OL_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIC_OL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHIC_OM_start                   : std_logic;
  signal AS_L2PHIC_OM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHIC_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHIC_OM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHIC_OM_wea          : t_AS_51_1b;
  signal AS_L2PHIC_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHIC_OM_din         : t_AS_51_DATA;
  signal AS_L2PHIC_OM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHIC_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHIC_OM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHIC_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHID_BM_start                   : std_logic;
  signal AS_L2PHID_BM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHID_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHID_BM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHID_BM_wea          : t_AS_51_1b;
  signal AS_L2PHID_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHID_BM_din         : t_AS_51_DATA;
  signal AS_L2PHID_BM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHID_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHID_BM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHID_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L2PHID_OM_start                   : std_logic;
  signal AS_L2PHID_OM_wea_delay          : t_AS_51_1b;
  signal AS_L2PHID_OM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L2PHID_OM_din_delay         : t_AS_51_DATA;
  signal AS_L2PHID_OM_wea          : t_AS_51_1b;
  signal AS_L2PHID_OM_writeaddr   : t_AS_51_ADDR;
  signal AS_L2PHID_OM_din         : t_AS_51_DATA;
  signal AS_L2PHID_OM_enb          : t_AS_51_1b := '1';
  signal AS_L2PHID_OM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L2PHID_OM_V_dout        : t_AS_51_DATA;
  signal AS_L2PHID_OM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L3PHIA_BM_start                   : std_logic;
  signal AS_L3PHIA_BM_wea_delay          : t_AS_51_1b;
  signal AS_L3PHIA_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L3PHIA_BM_din_delay         : t_AS_51_DATA;
  signal AS_L3PHIA_BM_wea          : t_AS_51_1b;
  signal AS_L3PHIA_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L3PHIA_BM_din         : t_AS_51_DATA;
  signal AS_L3PHIA_BM_enb          : t_AS_51_1b := '1';
  signal AS_L3PHIA_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L3PHIA_BM_V_dout        : t_AS_51_DATA;
  signal AS_L3PHIA_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L3PHIB_BM_start                   : std_logic;
  signal AS_L3PHIB_BM_wea_delay          : t_AS_51_1b;
  signal AS_L3PHIB_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L3PHIB_BM_din_delay         : t_AS_51_DATA;
  signal AS_L3PHIB_BM_wea          : t_AS_51_1b;
  signal AS_L3PHIB_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L3PHIB_BM_din         : t_AS_51_DATA;
  signal AS_L3PHIB_BM_enb          : t_AS_51_1b := '1';
  signal AS_L3PHIB_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L3PHIB_BM_V_dout        : t_AS_51_DATA;
  signal AS_L3PHIB_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L3PHIB_BR_start                   : std_logic;
  signal AS_L3PHIB_BR_wea_delay          : t_AS_51_1b;
  signal AS_L3PHIB_BR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L3PHIB_BR_din_delay         : t_AS_51_DATA;
  signal AS_L3PHIB_BR_wea          : t_AS_51_1b;
  signal AS_L3PHIB_BR_writeaddr   : t_AS_51_ADDR;
  signal AS_L3PHIB_BR_din         : t_AS_51_DATA;
  signal AS_L3PHIB_BR_enb          : t_AS_51_1b := '1';
  signal AS_L3PHIB_BR_V_readaddr    : t_AS_51_ADDR;
  signal AS_L3PHIB_BR_V_dout        : t_AS_51_DATA;
  signal AS_L3PHIB_BR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L3PHIC_BL_start                   : std_logic;
  signal AS_L3PHIC_BL_wea_delay          : t_AS_51_1b;
  signal AS_L3PHIC_BL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L3PHIC_BL_din_delay         : t_AS_51_DATA;
  signal AS_L3PHIC_BL_wea          : t_AS_51_1b;
  signal AS_L3PHIC_BL_writeaddr   : t_AS_51_ADDR;
  signal AS_L3PHIC_BL_din         : t_AS_51_DATA;
  signal AS_L3PHIC_BL_enb          : t_AS_51_1b := '1';
  signal AS_L3PHIC_BL_V_readaddr    : t_AS_51_ADDR;
  signal AS_L3PHIC_BL_V_dout        : t_AS_51_DATA;
  signal AS_L3PHIC_BL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L3PHIC_BM_start                   : std_logic;
  signal AS_L3PHIC_BM_wea_delay          : t_AS_51_1b;
  signal AS_L3PHIC_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L3PHIC_BM_din_delay         : t_AS_51_DATA;
  signal AS_L3PHIC_BM_wea          : t_AS_51_1b;
  signal AS_L3PHIC_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L3PHIC_BM_din         : t_AS_51_DATA;
  signal AS_L3PHIC_BM_enb          : t_AS_51_1b := '1';
  signal AS_L3PHIC_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L3PHIC_BM_V_dout        : t_AS_51_DATA;
  signal AS_L3PHIC_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L3PHID_BM_start                   : std_logic;
  signal AS_L3PHID_BM_wea_delay          : t_AS_51_1b;
  signal AS_L3PHID_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L3PHID_BM_din_delay         : t_AS_51_DATA;
  signal AS_L3PHID_BM_wea          : t_AS_51_1b;
  signal AS_L3PHID_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L3PHID_BM_din         : t_AS_51_DATA;
  signal AS_L3PHID_BM_enb          : t_AS_51_1b := '1';
  signal AS_L3PHID_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L3PHID_BM_V_dout        : t_AS_51_DATA;
  signal AS_L3PHID_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L5PHIA_BM_start                   : std_logic;
  signal AS_L5PHIA_BM_wea_delay          : t_AS_51_1b;
  signal AS_L5PHIA_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L5PHIA_BM_din_delay         : t_AS_51_DATA;
  signal AS_L5PHIA_BM_wea          : t_AS_51_1b;
  signal AS_L5PHIA_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L5PHIA_BM_din         : t_AS_51_DATA;
  signal AS_L5PHIA_BM_enb          : t_AS_51_1b := '1';
  signal AS_L5PHIA_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L5PHIA_BM_V_dout        : t_AS_51_DATA;
  signal AS_L5PHIA_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L5PHIB_BM_start                   : std_logic;
  signal AS_L5PHIB_BM_wea_delay          : t_AS_51_1b;
  signal AS_L5PHIB_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L5PHIB_BM_din_delay         : t_AS_51_DATA;
  signal AS_L5PHIB_BM_wea          : t_AS_51_1b;
  signal AS_L5PHIB_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L5PHIB_BM_din         : t_AS_51_DATA;
  signal AS_L5PHIB_BM_enb          : t_AS_51_1b := '1';
  signal AS_L5PHIB_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L5PHIB_BM_V_dout        : t_AS_51_DATA;
  signal AS_L5PHIB_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L5PHIB_BR_start                   : std_logic;
  signal AS_L5PHIB_BR_wea_delay          : t_AS_51_1b;
  signal AS_L5PHIB_BR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L5PHIB_BR_din_delay         : t_AS_51_DATA;
  signal AS_L5PHIB_BR_wea          : t_AS_51_1b;
  signal AS_L5PHIB_BR_writeaddr   : t_AS_51_ADDR;
  signal AS_L5PHIB_BR_din         : t_AS_51_DATA;
  signal AS_L5PHIB_BR_enb          : t_AS_51_1b := '1';
  signal AS_L5PHIB_BR_V_readaddr    : t_AS_51_ADDR;
  signal AS_L5PHIB_BR_V_dout        : t_AS_51_DATA;
  signal AS_L5PHIB_BR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L5PHIC_BL_start                   : std_logic;
  signal AS_L5PHIC_BL_wea_delay          : t_AS_51_1b;
  signal AS_L5PHIC_BL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L5PHIC_BL_din_delay         : t_AS_51_DATA;
  signal AS_L5PHIC_BL_wea          : t_AS_51_1b;
  signal AS_L5PHIC_BL_writeaddr   : t_AS_51_ADDR;
  signal AS_L5PHIC_BL_din         : t_AS_51_DATA;
  signal AS_L5PHIC_BL_enb          : t_AS_51_1b := '1';
  signal AS_L5PHIC_BL_V_readaddr    : t_AS_51_ADDR;
  signal AS_L5PHIC_BL_V_dout        : t_AS_51_DATA;
  signal AS_L5PHIC_BL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L5PHIC_BM_start                   : std_logic;
  signal AS_L5PHIC_BM_wea_delay          : t_AS_51_1b;
  signal AS_L5PHIC_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L5PHIC_BM_din_delay         : t_AS_51_DATA;
  signal AS_L5PHIC_BM_wea          : t_AS_51_1b;
  signal AS_L5PHIC_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L5PHIC_BM_din         : t_AS_51_DATA;
  signal AS_L5PHIC_BM_enb          : t_AS_51_1b := '1';
  signal AS_L5PHIC_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L5PHIC_BM_V_dout        : t_AS_51_DATA;
  signal AS_L5PHIC_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_L5PHID_BM_start                   : std_logic;
  signal AS_L5PHID_BM_wea_delay          : t_AS_51_1b;
  signal AS_L5PHID_BM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_L5PHID_BM_din_delay         : t_AS_51_DATA;
  signal AS_L5PHID_BM_wea          : t_AS_51_1b;
  signal AS_L5PHID_BM_writeaddr   : t_AS_51_ADDR;
  signal AS_L5PHID_BM_din         : t_AS_51_DATA;
  signal AS_L5PHID_BM_enb          : t_AS_51_1b := '1';
  signal AS_L5PHID_BM_V_readaddr    : t_AS_51_ADDR;
  signal AS_L5PHID_BM_V_dout        : t_AS_51_DATA;
  signal AS_L5PHID_BM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D1PHIA_DM_start                   : std_logic;
  signal AS_D1PHIA_DM_wea_delay          : t_AS_51_1b;
  signal AS_D1PHIA_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D1PHIA_DM_din_delay         : t_AS_51_DATA;
  signal AS_D1PHIA_DM_wea          : t_AS_51_1b;
  signal AS_D1PHIA_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D1PHIA_DM_din         : t_AS_51_DATA;
  signal AS_D1PHIA_DM_enb          : t_AS_51_1b := '1';
  signal AS_D1PHIA_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D1PHIA_DM_V_dout        : t_AS_51_DATA;
  signal AS_D1PHIA_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D1PHIB_DM_start                   : std_logic;
  signal AS_D1PHIB_DM_wea_delay          : t_AS_51_1b;
  signal AS_D1PHIB_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D1PHIB_DM_din_delay         : t_AS_51_DATA;
  signal AS_D1PHIB_DM_wea          : t_AS_51_1b;
  signal AS_D1PHIB_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D1PHIB_DM_din         : t_AS_51_DATA;
  signal AS_D1PHIB_DM_enb          : t_AS_51_1b := '1';
  signal AS_D1PHIB_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D1PHIB_DM_V_dout        : t_AS_51_DATA;
  signal AS_D1PHIB_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D1PHIB_DR_start                   : std_logic;
  signal AS_D1PHIB_DR_wea_delay          : t_AS_51_1b;
  signal AS_D1PHIB_DR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D1PHIB_DR_din_delay         : t_AS_51_DATA;
  signal AS_D1PHIB_DR_wea          : t_AS_51_1b;
  signal AS_D1PHIB_DR_writeaddr   : t_AS_51_ADDR;
  signal AS_D1PHIB_DR_din         : t_AS_51_DATA;
  signal AS_D1PHIB_DR_enb          : t_AS_51_1b := '1';
  signal AS_D1PHIB_DR_V_readaddr    : t_AS_51_ADDR;
  signal AS_D1PHIB_DR_V_dout        : t_AS_51_DATA;
  signal AS_D1PHIB_DR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D1PHIC_DL_start                   : std_logic;
  signal AS_D1PHIC_DL_wea_delay          : t_AS_51_1b;
  signal AS_D1PHIC_DL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D1PHIC_DL_din_delay         : t_AS_51_DATA;
  signal AS_D1PHIC_DL_wea          : t_AS_51_1b;
  signal AS_D1PHIC_DL_writeaddr   : t_AS_51_ADDR;
  signal AS_D1PHIC_DL_din         : t_AS_51_DATA;
  signal AS_D1PHIC_DL_enb          : t_AS_51_1b := '1';
  signal AS_D1PHIC_DL_V_readaddr    : t_AS_51_ADDR;
  signal AS_D1PHIC_DL_V_dout        : t_AS_51_DATA;
  signal AS_D1PHIC_DL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D1PHIC_DM_start                   : std_logic;
  signal AS_D1PHIC_DM_wea_delay          : t_AS_51_1b;
  signal AS_D1PHIC_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D1PHIC_DM_din_delay         : t_AS_51_DATA;
  signal AS_D1PHIC_DM_wea          : t_AS_51_1b;
  signal AS_D1PHIC_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D1PHIC_DM_din         : t_AS_51_DATA;
  signal AS_D1PHIC_DM_enb          : t_AS_51_1b := '1';
  signal AS_D1PHIC_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D1PHIC_DM_V_dout        : t_AS_51_DATA;
  signal AS_D1PHIC_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D1PHID_DM_start                   : std_logic;
  signal AS_D1PHID_DM_wea_delay          : t_AS_51_1b;
  signal AS_D1PHID_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D1PHID_DM_din_delay         : t_AS_51_DATA;
  signal AS_D1PHID_DM_wea          : t_AS_51_1b;
  signal AS_D1PHID_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D1PHID_DM_din         : t_AS_51_DATA;
  signal AS_D1PHID_DM_enb          : t_AS_51_1b := '1';
  signal AS_D1PHID_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D1PHID_DM_V_dout        : t_AS_51_DATA;
  signal AS_D1PHID_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D3PHIA_DM_start                   : std_logic;
  signal AS_D3PHIA_DM_wea_delay          : t_AS_51_1b;
  signal AS_D3PHIA_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D3PHIA_DM_din_delay         : t_AS_51_DATA;
  signal AS_D3PHIA_DM_wea          : t_AS_51_1b;
  signal AS_D3PHIA_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D3PHIA_DM_din         : t_AS_51_DATA;
  signal AS_D3PHIA_DM_enb          : t_AS_51_1b := '1';
  signal AS_D3PHIA_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D3PHIA_DM_V_dout        : t_AS_51_DATA;
  signal AS_D3PHIA_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D3PHIB_DM_start                   : std_logic;
  signal AS_D3PHIB_DM_wea_delay          : t_AS_51_1b;
  signal AS_D3PHIB_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D3PHIB_DM_din_delay         : t_AS_51_DATA;
  signal AS_D3PHIB_DM_wea          : t_AS_51_1b;
  signal AS_D3PHIB_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D3PHIB_DM_din         : t_AS_51_DATA;
  signal AS_D3PHIB_DM_enb          : t_AS_51_1b := '1';
  signal AS_D3PHIB_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D3PHIB_DM_V_dout        : t_AS_51_DATA;
  signal AS_D3PHIB_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D3PHIB_DR_start                   : std_logic;
  signal AS_D3PHIB_DR_wea_delay          : t_AS_51_1b;
  signal AS_D3PHIB_DR_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D3PHIB_DR_din_delay         : t_AS_51_DATA;
  signal AS_D3PHIB_DR_wea          : t_AS_51_1b;
  signal AS_D3PHIB_DR_writeaddr   : t_AS_51_ADDR;
  signal AS_D3PHIB_DR_din         : t_AS_51_DATA;
  signal AS_D3PHIB_DR_enb          : t_AS_51_1b := '1';
  signal AS_D3PHIB_DR_V_readaddr    : t_AS_51_ADDR;
  signal AS_D3PHIB_DR_V_dout        : t_AS_51_DATA;
  signal AS_D3PHIB_DR_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D3PHIC_DL_start                   : std_logic;
  signal AS_D3PHIC_DL_wea_delay          : t_AS_51_1b;
  signal AS_D3PHIC_DL_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D3PHIC_DL_din_delay         : t_AS_51_DATA;
  signal AS_D3PHIC_DL_wea          : t_AS_51_1b;
  signal AS_D3PHIC_DL_writeaddr   : t_AS_51_ADDR;
  signal AS_D3PHIC_DL_din         : t_AS_51_DATA;
  signal AS_D3PHIC_DL_enb          : t_AS_51_1b := '1';
  signal AS_D3PHIC_DL_V_readaddr    : t_AS_51_ADDR;
  signal AS_D3PHIC_DL_V_dout        : t_AS_51_DATA;
  signal AS_D3PHIC_DL_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D3PHIC_DM_start                   : std_logic;
  signal AS_D3PHIC_DM_wea_delay          : t_AS_51_1b;
  signal AS_D3PHIC_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D3PHIC_DM_din_delay         : t_AS_51_DATA;
  signal AS_D3PHIC_DM_wea          : t_AS_51_1b;
  signal AS_D3PHIC_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D3PHIC_DM_din         : t_AS_51_DATA;
  signal AS_D3PHIC_DM_enb          : t_AS_51_1b := '1';
  signal AS_D3PHIC_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D3PHIC_DM_V_dout        : t_AS_51_DATA;
  signal AS_D3PHIC_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal AS_D3PHID_DM_start                   : std_logic;
  signal AS_D3PHID_DM_wea_delay          : t_AS_51_1b;
  signal AS_D3PHID_DM_writeaddr_delay   : t_AS_51_ADDR;
  signal AS_D3PHID_DM_din_delay         : t_AS_51_DATA;
  signal AS_D3PHID_DM_wea          : t_AS_51_1b;
  signal AS_D3PHID_DM_writeaddr   : t_AS_51_ADDR;
  signal AS_D3PHID_DM_din         : t_AS_51_DATA;
  signal AS_D3PHID_DM_enb          : t_AS_51_1b := '1';
  signal AS_D3PHID_DM_V_readaddr    : t_AS_51_ADDR;
  signal AS_D3PHID_DM_V_dout        : t_AS_51_DATA;
  signal AS_D3PHID_DM_AV_dout_nent  : t_AS_51_NENT; -- (#page)
  signal VMSTE_L2PHIAn1_start                   : std_logic;
  signal VMSTE_L2PHIAn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIAn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIAn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIAn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIAn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIAn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIAn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIAn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIAn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIAn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIAn1_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIAn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIAn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIAn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIAn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIAn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIAn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn2_start                   : std_logic;
  signal VMSTE_L2PHIAn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIAn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIAn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIAn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIAn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIAn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIAn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIAn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIAn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIAn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIAn2_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIAn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIAn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIAn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIAn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIAn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIAn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn3_start                   : std_logic;
  signal VMSTE_L2PHIAn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIAn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIAn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIAn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIAn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIAn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIAn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIAn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIAn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIAn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIAn3_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIAn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIAn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIAn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIAn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIAn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIAn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIAn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn1_start                   : std_logic;
  signal VMSTE_L2PHIBn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIBn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIBn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIBn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIBn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIBn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIBn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIBn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIBn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIBn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIBn1_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIBn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIBn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIBn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIBn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIBn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIBn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn2_start                   : std_logic;
  signal VMSTE_L2PHIBn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIBn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIBn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIBn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIBn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIBn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIBn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIBn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIBn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIBn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIBn2_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIBn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIBn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIBn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIBn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIBn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIBn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn3_start                   : std_logic;
  signal VMSTE_L2PHIBn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIBn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIBn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIBn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIBn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIBn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIBn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIBn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIBn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIBn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIBn3_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIBn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIBn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIBn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIBn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIBn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIBn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIBn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn1_start                   : std_logic;
  signal VMSTE_L2PHICn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHICn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHICn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHICn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHICn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHICn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHICn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHICn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHICn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHICn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHICn1_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHICn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHICn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHICn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHICn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHICn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHICn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn2_start                   : std_logic;
  signal VMSTE_L2PHICn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHICn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHICn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHICn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHICn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHICn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHICn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHICn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHICn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHICn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHICn2_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHICn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHICn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHICn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHICn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHICn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHICn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn3_start                   : std_logic;
  signal VMSTE_L2PHICn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHICn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHICn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHICn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHICn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHICn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHICn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHICn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHICn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHICn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHICn3_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHICn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHICn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHICn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHICn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHICn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHICn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHICn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn1_start                   : std_logic;
  signal VMSTE_L2PHIDn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIDn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIDn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIDn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIDn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIDn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIDn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIDn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIDn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIDn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIDn1_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIDn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIDn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIDn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIDn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIDn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIDn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn2_start                   : std_logic;
  signal VMSTE_L2PHIDn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIDn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIDn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIDn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIDn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIDn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIDn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIDn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIDn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIDn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIDn2_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIDn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIDn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIDn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIDn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIDn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIDn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn3_start                   : std_logic;
  signal VMSTE_L2PHIDn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIDn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIDn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L2PHIDn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_L2PHIDn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L2PHIDn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L2PHIDn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L2PHIDn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L2PHIDn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L2PHIDn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L2PHIDn3_V_datatmp : t_VMSTE_16_DATA_5;
  signal VMSTE_L2PHIDn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L2PHIDn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIDn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIDn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L2PHIDn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L2PHIDn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L2PHIDn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L3PHIIn1_start                   : std_logic;
  signal VMSTE_L3PHIIn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L3PHIIn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHIIn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHIIn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L3PHIIn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHIIn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHIIn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L3PHIIn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L3PHIIn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L3PHIIn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L3PHIIn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L3PHIIn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L3PHIIn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L3PHIIn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_L3PHIIn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L3PHIIn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHIIn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHIIn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L3PHIIn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHIIn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHIIn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L3PHIJn1_start                   : std_logic;
  signal VMSTE_L3PHIJn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L3PHIJn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHIJn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHIJn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L3PHIJn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHIJn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHIJn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L3PHIJn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L3PHIJn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L3PHIJn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L3PHIJn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L3PHIJn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L3PHIJn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L3PHIJn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_L3PHIJn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L3PHIJn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHIJn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHIJn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L3PHIJn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHIJn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHIJn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L3PHIKn1_start                   : std_logic;
  signal VMSTE_L3PHIKn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L3PHIKn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHIKn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHIKn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L3PHIKn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHIKn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHIKn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L3PHIKn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L3PHIKn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L3PHIKn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L3PHIKn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L3PHIKn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L3PHIKn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L3PHIKn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_L3PHIKn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L3PHIKn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHIKn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHIKn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L3PHIKn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHIKn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHIKn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L3PHILn1_start                   : std_logic;
  signal VMSTE_L3PHILn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_L3PHILn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHILn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHILn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_L3PHILn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_L3PHILn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_L3PHILn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_L3PHILn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_L3PHILn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_L3PHILn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_L3PHILn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_L3PHILn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_L3PHILn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_L3PHILn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_L3PHILn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_L3PHILn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHILn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHILn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_L3PHILn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_L3PHILn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_L3PHILn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D2PHIAn1_start                   : std_logic;
  signal VMSTE_D2PHIAn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D2PHIAn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHIAn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHIAn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D2PHIAn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHIAn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHIAn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D2PHIAn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D2PHIAn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D2PHIAn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D2PHIAn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D2PHIAn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D2PHIAn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D2PHIAn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D2PHIAn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D2PHIAn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHIAn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHIAn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D2PHIAn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHIAn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHIAn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D2PHIBn1_start                   : std_logic;
  signal VMSTE_D2PHIBn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D2PHIBn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHIBn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHIBn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D2PHIBn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHIBn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHIBn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D2PHIBn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D2PHIBn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D2PHIBn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D2PHIBn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D2PHIBn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D2PHIBn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D2PHIBn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D2PHIBn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D2PHIBn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHIBn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHIBn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D2PHIBn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHIBn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHIBn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D2PHICn1_start                   : std_logic;
  signal VMSTE_D2PHICn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D2PHICn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHICn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHICn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D2PHICn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHICn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHICn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D2PHICn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D2PHICn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D2PHICn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D2PHICn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D2PHICn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D2PHICn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D2PHICn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D2PHICn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D2PHICn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHICn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHICn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D2PHICn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHICn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHICn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D2PHIDn1_start                   : std_logic;
  signal VMSTE_D2PHIDn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D2PHIDn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHIDn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHIDn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D2PHIDn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D2PHIDn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D2PHIDn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D2PHIDn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D2PHIDn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D2PHIDn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D2PHIDn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D2PHIDn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D2PHIDn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D2PHIDn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D2PHIDn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D2PHIDn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHIDn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHIDn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D2PHIDn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D2PHIDn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D2PHIDn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D4PHIAn1_start                   : std_logic;
  signal VMSTE_D4PHIAn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D4PHIAn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHIAn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHIAn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D4PHIAn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHIAn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHIAn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D4PHIAn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D4PHIAn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D4PHIAn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D4PHIAn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D4PHIAn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D4PHIAn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D4PHIAn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D4PHIAn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D4PHIAn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHIAn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHIAn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D4PHIAn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHIAn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHIAn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D4PHIBn1_start                   : std_logic;
  signal VMSTE_D4PHIBn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D4PHIBn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHIBn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHIBn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D4PHIBn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHIBn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHIBn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D4PHIBn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D4PHIBn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D4PHIBn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D4PHIBn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D4PHIBn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D4PHIBn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D4PHIBn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D4PHIBn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D4PHIBn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHIBn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHIBn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D4PHIBn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHIBn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHIBn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D4PHICn1_start                   : std_logic;
  signal VMSTE_D4PHICn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D4PHICn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHICn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHICn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D4PHICn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHICn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHICn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D4PHICn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D4PHICn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D4PHICn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D4PHICn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D4PHICn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D4PHICn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D4PHICn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D4PHICn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D4PHICn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHICn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHICn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D4PHICn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHICn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHICn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D4PHIDn1_start                   : std_logic;
  signal VMSTE_D4PHIDn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D4PHIDn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHIDn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHIDn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D4PHIDn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D4PHIDn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D4PHIDn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D4PHIDn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D4PHIDn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D4PHIDn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D4PHIDn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D4PHIDn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D4PHIDn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D4PHIDn1_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D4PHIDn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D4PHIDn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHIDn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHIDn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D4PHIDn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D4PHIDn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D4PHIDn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn1_start                   : std_logic;
  signal VMSTE_D1PHIXn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIXn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIXn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIXn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIXn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIXn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIXn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIXn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIXn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIXn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIXn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIXn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIXn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIXn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIXn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIXn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIXn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn2_start                   : std_logic;
  signal VMSTE_D1PHIXn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIXn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIXn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIXn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIXn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIXn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIXn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIXn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIXn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIXn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIXn2_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIXn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIXn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIXn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIXn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIXn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIXn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn1_start                   : std_logic;
  signal VMSTE_D1PHIYn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIYn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIYn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIYn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIYn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIYn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIYn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIYn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIYn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIYn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIYn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIYn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIYn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIYn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIYn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIYn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIYn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn2_start                   : std_logic;
  signal VMSTE_D1PHIYn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIYn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIYn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIYn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIYn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIYn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIYn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIYn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIYn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIYn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIYn2_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIYn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIYn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIYn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIYn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIYn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIYn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn1_start                   : std_logic;
  signal VMSTE_D1PHIZn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIZn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIZn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIZn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIZn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIZn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIZn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIZn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIZn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIZn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIZn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIZn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIZn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIZn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIZn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIZn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIZn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn2_start                   : std_logic;
  signal VMSTE_D1PHIZn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIZn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIZn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIZn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIZn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIZn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIZn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIZn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIZn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIZn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIZn2_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIZn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIZn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIZn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIZn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIZn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIZn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn1_start                   : std_logic;
  signal VMSTE_D1PHIWn1_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn1_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIWn1_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIWn1_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn1_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIWn1_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIWn1_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIWn1_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIWn1_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIWn1_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIWn1_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn1_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIWn1_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIWn1_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIWn1_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIWn1_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIWn1_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIWn1_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn1_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIWn1_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIWn1_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn2_start                   : std_logic;
  signal VMSTE_D1PHIWn2_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn2_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIWn2_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIWn2_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn2_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIWn2_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIWn2_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIWn2_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIWn2_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIWn2_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIWn2_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn2_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIWn2_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIWn2_V_datatmp : t_VMSTE_16_DATA_3;
  signal VMSTE_D1PHIWn2_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIWn2_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIWn2_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIWn2_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn2_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIWn2_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIWn2_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn3_start                   : std_logic;
  signal VMSTE_D1PHIXn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIXn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIXn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIXn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIXn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIXn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIXn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIXn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIXn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIXn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIXn3_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D1PHIXn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIXn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIXn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIXn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIXn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIXn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIXn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn3_start                   : std_logic;
  signal VMSTE_D1PHIYn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIYn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIYn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIYn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIYn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIYn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIYn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIYn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIYn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIYn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIYn3_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D1PHIYn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIYn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIYn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIYn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIYn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIYn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIYn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn3_start                   : std_logic;
  signal VMSTE_D1PHIZn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIZn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIZn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIZn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIZn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIZn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIZn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIZn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIZn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIZn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIZn3_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D1PHIZn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIZn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIZn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIZn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIZn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIZn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIZn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn3_start                   : std_logic;
  signal VMSTE_D1PHIWn3_wea_delay          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn3_writeaddr_delay   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIWn3_din_delay         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIWn3_wea          : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn3_writeaddr   : t_VMSTE_16_ADDR;
  signal VMSTE_D1PHIWn3_din         : t_VMSTE_16_DATA;
  signal VMSTE_D1PHIWn3_A_enb         : t_VMSTE_16_A1b;
  signal VMSTE_D1PHIWn3_AV_readaddr   : t_VMSTE_16_AADDR;
  signal VMSTE_D1PHIWn3_AV_dout       : t_VMSTE_16_ADATA;
  signal VMSTE_D1PHIWn3_AV_dout_mask : t_VMSTE_16_MASK; -- (#page)(#bin)
  signal VMSTE_D1PHIWn3_enb_nent         : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn3_V_addr_nent   : t_VMSTE_16_NENTADDR;
  signal VMSTE_D1PHIWn3_AV_dout_nent : t_VMSTE_16_NENT; -- (#page)(#bin)
  signal VMSTE_D1PHIWn3_V_datatmp : t_VMSTE_16_DATA_2;
  signal VMSTE_D1PHIWn3_V_masktmp : t_VMSTE_16_MASK_2;
  signal VMSTE_D1PHIWn3_V_addr_binmaskA   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIWn3_V_binmaskA   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIWn3_enb_binmaskA   : t_VMSTE_16_1b;
  signal VMSTE_D1PHIWn3_V_addr_binmaskB   : t_VMSTE_16_ADDRBINMASK;
  signal VMSTE_D1PHIWn3_V_binmaskB   : t_VMSTE_16_BINMASK;
  signal VMSTE_D1PHIWn3_enb_binmaskB   : t_VMSTE_16_1b;
  signal VMSTE_L4PHIAn1_start                   : std_logic;
  signal VMSTE_L4PHIAn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L4PHIAn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHIAn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHIAn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L4PHIAn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHIAn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHIAn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L4PHIAn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L4PHIAn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L4PHIAn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L4PHIAn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L4PHIAn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L4PHIAn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L4PHIAn1_V_datatmp : t_VMSTE_17_DATA_5;
  signal VMSTE_L4PHIAn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L4PHIAn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHIAn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHIAn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L4PHIAn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHIAn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHIAn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal VMSTE_L4PHIBn1_start                   : std_logic;
  signal VMSTE_L4PHIBn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L4PHIBn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHIBn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHIBn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L4PHIBn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHIBn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHIBn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L4PHIBn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L4PHIBn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L4PHIBn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L4PHIBn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L4PHIBn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L4PHIBn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L4PHIBn1_V_datatmp : t_VMSTE_17_DATA_5;
  signal VMSTE_L4PHIBn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L4PHIBn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHIBn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHIBn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L4PHIBn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHIBn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHIBn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal VMSTE_L4PHICn1_start                   : std_logic;
  signal VMSTE_L4PHICn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L4PHICn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHICn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHICn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L4PHICn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHICn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHICn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L4PHICn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L4PHICn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L4PHICn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L4PHICn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L4PHICn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L4PHICn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L4PHICn1_V_datatmp : t_VMSTE_17_DATA_5;
  signal VMSTE_L4PHICn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L4PHICn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHICn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHICn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L4PHICn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHICn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHICn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal VMSTE_L4PHIDn1_start                   : std_logic;
  signal VMSTE_L4PHIDn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L4PHIDn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHIDn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHIDn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L4PHIDn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L4PHIDn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L4PHIDn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L4PHIDn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L4PHIDn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L4PHIDn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L4PHIDn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L4PHIDn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L4PHIDn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L4PHIDn1_V_datatmp : t_VMSTE_17_DATA_5;
  signal VMSTE_L4PHIDn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L4PHIDn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHIDn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHIDn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L4PHIDn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L4PHIDn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L4PHIDn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal VMSTE_L6PHIAn1_start                   : std_logic;
  signal VMSTE_L6PHIAn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L6PHIAn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHIAn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHIAn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L6PHIAn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHIAn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHIAn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L6PHIAn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L6PHIAn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L6PHIAn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L6PHIAn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L6PHIAn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L6PHIAn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L6PHIAn1_V_datatmp : t_VMSTE_17_DATA_3;
  signal VMSTE_L6PHIAn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L6PHIAn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHIAn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHIAn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L6PHIAn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHIAn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHIAn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal VMSTE_L6PHIBn1_start                   : std_logic;
  signal VMSTE_L6PHIBn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L6PHIBn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHIBn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHIBn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L6PHIBn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHIBn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHIBn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L6PHIBn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L6PHIBn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L6PHIBn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L6PHIBn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L6PHIBn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L6PHIBn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L6PHIBn1_V_datatmp : t_VMSTE_17_DATA_3;
  signal VMSTE_L6PHIBn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L6PHIBn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHIBn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHIBn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L6PHIBn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHIBn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHIBn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal VMSTE_L6PHICn1_start                   : std_logic;
  signal VMSTE_L6PHICn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L6PHICn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHICn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHICn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L6PHICn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHICn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHICn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L6PHICn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L6PHICn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L6PHICn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L6PHICn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L6PHICn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L6PHICn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L6PHICn1_V_datatmp : t_VMSTE_17_DATA_3;
  signal VMSTE_L6PHICn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L6PHICn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHICn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHICn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L6PHICn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHICn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHICn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal VMSTE_L6PHIDn1_start                   : std_logic;
  signal VMSTE_L6PHIDn1_wea_delay          : t_VMSTE_17_1b;
  signal VMSTE_L6PHIDn1_writeaddr_delay   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHIDn1_din_delay         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHIDn1_wea          : t_VMSTE_17_1b;
  signal VMSTE_L6PHIDn1_writeaddr   : t_VMSTE_17_ADDR;
  signal VMSTE_L6PHIDn1_din         : t_VMSTE_17_DATA;
  signal VMSTE_L6PHIDn1_A_enb         : t_VMSTE_17_A1b;
  signal VMSTE_L6PHIDn1_AV_readaddr   : t_VMSTE_17_AADDR;
  signal VMSTE_L6PHIDn1_AV_dout       : t_VMSTE_17_ADATA;
  signal VMSTE_L6PHIDn1_AV_dout_mask : t_VMSTE_17_MASK; -- (#page)(#bin)
  signal VMSTE_L6PHIDn1_enb_nent         : t_VMSTE_17_1b;
  signal VMSTE_L6PHIDn1_V_addr_nent   : t_VMSTE_17_NENTADDR;
  signal VMSTE_L6PHIDn1_AV_dout_nent : t_VMSTE_17_NENT; -- (#page)(#bin)
  signal VMSTE_L6PHIDn1_V_datatmp : t_VMSTE_17_DATA_3;
  signal VMSTE_L6PHIDn1_V_masktmp : t_VMSTE_17_MASK_2;
  signal VMSTE_L6PHIDn1_V_addr_binmaskA   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHIDn1_V_binmaskA   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHIDn1_enb_binmaskA   : t_VMSTE_17_1b;
  signal VMSTE_L6PHIDn1_V_addr_binmaskB   : t_VMSTE_17_ADDRBINMASK;
  signal VMSTE_L6PHIDn1_V_binmaskB   : t_VMSTE_17_BINMASK;
  signal VMSTE_L6PHIDn1_enb_binmaskB   : t_VMSTE_17_1b;
  signal TPAR_L1L2A_start                   : std_logic;
  signal TPAR_L1L2A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2A_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2A_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2B_start                   : std_logic;
  signal TPAR_L1L2B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2B_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2B_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2C_start                   : std_logic;
  signal TPAR_L1L2C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2C_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2C_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2D_start                   : std_logic;
  signal TPAR_L1L2D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2D_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2D_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2E_start                   : std_logic;
  signal TPAR_L1L2E_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2E_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2E_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2E_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2E_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2E_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2E_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2E_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2E_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2E_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2E_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2F_start                   : std_logic;
  signal TPAR_L1L2F_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2F_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2F_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2F_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2F_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2F_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2F_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2F_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2F_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2F_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2F_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2G_start                   : std_logic;
  signal TPAR_L1L2G_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2G_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2G_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2G_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2G_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2G_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2G_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2G_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2G_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2G_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2G_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2H_start                   : std_logic;
  signal TPAR_L1L2H_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2H_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2H_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2H_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2H_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2H_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2H_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2H_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2H_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2H_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2H_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2I_start                   : std_logic;
  signal TPAR_L1L2I_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2I_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2I_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2I_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2I_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2I_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2I_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2I_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2I_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2I_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2I_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2J_start                   : std_logic;
  signal TPAR_L1L2J_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2J_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2J_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2J_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2J_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2J_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2J_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2J_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2J_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2J_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2J_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2K_start                   : std_logic;
  signal TPAR_L1L2K_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2K_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2K_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2K_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2K_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2K_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2K_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2K_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2K_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2K_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2K_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1L2L_start                   : std_logic;
  signal TPAR_L1L2L_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1L2L_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1L2L_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1L2L_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1L2L_wea          : t_TPAR_73_1b;
  signal TPAR_L1L2L_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1L2L_din         : t_TPAR_73_DATA;
  signal TPAR_L1L2L_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1L2L_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1L2L_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1L2L_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2L3A_start                   : std_logic;
  signal TPAR_L2L3A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2L3A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2L3A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2L3A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2L3A_wea          : t_TPAR_73_1b;
  signal TPAR_L2L3A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2L3A_din         : t_TPAR_73_DATA;
  signal TPAR_L2L3A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2L3A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2L3A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2L3A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2L3B_start                   : std_logic;
  signal TPAR_L2L3B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2L3B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2L3B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2L3B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2L3B_wea          : t_TPAR_73_1b;
  signal TPAR_L2L3B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2L3B_din         : t_TPAR_73_DATA;
  signal TPAR_L2L3B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2L3B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2L3B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2L3B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2L3C_start                   : std_logic;
  signal TPAR_L2L3C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2L3C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2L3C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2L3C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2L3C_wea          : t_TPAR_73_1b;
  signal TPAR_L2L3C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2L3C_din         : t_TPAR_73_DATA;
  signal TPAR_L2L3C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2L3C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2L3C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2L3C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2L3D_start                   : std_logic;
  signal TPAR_L2L3D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2L3D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2L3D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2L3D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2L3D_wea          : t_TPAR_73_1b;
  signal TPAR_L2L3D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2L3D_din         : t_TPAR_73_DATA;
  signal TPAR_L2L3D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2L3D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2L3D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2L3D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L3L4A_start                   : std_logic;
  signal TPAR_L3L4A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L3L4A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L3L4A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L3L4A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L3L4A_wea          : t_TPAR_73_1b;
  signal TPAR_L3L4A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L3L4A_din         : t_TPAR_73_DATA;
  signal TPAR_L3L4A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L3L4A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L3L4A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L3L4A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L3L4B_start                   : std_logic;
  signal TPAR_L3L4B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L3L4B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L3L4B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L3L4B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L3L4B_wea          : t_TPAR_73_1b;
  signal TPAR_L3L4B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L3L4B_din         : t_TPAR_73_DATA;
  signal TPAR_L3L4B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L3L4B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L3L4B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L3L4B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L3L4C_start                   : std_logic;
  signal TPAR_L3L4C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L3L4C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L3L4C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L3L4C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L3L4C_wea          : t_TPAR_73_1b;
  signal TPAR_L3L4C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L3L4C_din         : t_TPAR_73_DATA;
  signal TPAR_L3L4C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L3L4C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L3L4C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L3L4C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L3L4D_start                   : std_logic;
  signal TPAR_L3L4D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L3L4D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L3L4D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L3L4D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L3L4D_wea          : t_TPAR_73_1b;
  signal TPAR_L3L4D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L3L4D_din         : t_TPAR_73_DATA;
  signal TPAR_L3L4D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L3L4D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L3L4D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L3L4D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L5L6A_start                   : std_logic;
  signal TPAR_L5L6A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L5L6A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L5L6A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L5L6A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L5L6A_wea          : t_TPAR_73_1b;
  signal TPAR_L5L6A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L5L6A_din         : t_TPAR_73_DATA;
  signal TPAR_L5L6A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L5L6A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L5L6A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L5L6A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L5L6B_start                   : std_logic;
  signal TPAR_L5L6B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L5L6B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L5L6B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L5L6B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L5L6B_wea          : t_TPAR_73_1b;
  signal TPAR_L5L6B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L5L6B_din         : t_TPAR_73_DATA;
  signal TPAR_L5L6B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L5L6B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L5L6B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L5L6B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L5L6C_start                   : std_logic;
  signal TPAR_L5L6C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L5L6C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L5L6C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L5L6C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L5L6C_wea          : t_TPAR_73_1b;
  signal TPAR_L5L6C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L5L6C_din         : t_TPAR_73_DATA;
  signal TPAR_L5L6C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L5L6C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L5L6C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L5L6C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L5L6D_start                   : std_logic;
  signal TPAR_L5L6D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L5L6D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L5L6D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L5L6D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L5L6D_wea          : t_TPAR_73_1b;
  signal TPAR_L5L6D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L5L6D_din         : t_TPAR_73_DATA;
  signal TPAR_L5L6D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L5L6D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L5L6D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L5L6D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D1D2A_start                   : std_logic;
  signal TPAR_D1D2A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D1D2A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D1D2A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D1D2A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D1D2A_wea          : t_TPAR_73_1b;
  signal TPAR_D1D2A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D1D2A_din         : t_TPAR_73_DATA;
  signal TPAR_D1D2A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D1D2A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D1D2A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D1D2A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D1D2B_start                   : std_logic;
  signal TPAR_D1D2B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D1D2B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D1D2B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D1D2B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D1D2B_wea          : t_TPAR_73_1b;
  signal TPAR_D1D2B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D1D2B_din         : t_TPAR_73_DATA;
  signal TPAR_D1D2B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D1D2B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D1D2B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D1D2B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D1D2C_start                   : std_logic;
  signal TPAR_D1D2C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D1D2C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D1D2C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D1D2C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D1D2C_wea          : t_TPAR_73_1b;
  signal TPAR_D1D2C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D1D2C_din         : t_TPAR_73_DATA;
  signal TPAR_D1D2C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D1D2C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D1D2C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D1D2C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D1D2D_start                   : std_logic;
  signal TPAR_D1D2D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D1D2D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D1D2D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D1D2D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D1D2D_wea          : t_TPAR_73_1b;
  signal TPAR_D1D2D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D1D2D_din         : t_TPAR_73_DATA;
  signal TPAR_D1D2D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D1D2D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D1D2D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D1D2D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D3D4A_start                   : std_logic;
  signal TPAR_D3D4A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D3D4A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D3D4A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D3D4A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D3D4A_wea          : t_TPAR_73_1b;
  signal TPAR_D3D4A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D3D4A_din         : t_TPAR_73_DATA;
  signal TPAR_D3D4A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D3D4A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D3D4A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D3D4A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D3D4B_start                   : std_logic;
  signal TPAR_D3D4B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D3D4B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D3D4B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D3D4B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D3D4B_wea          : t_TPAR_73_1b;
  signal TPAR_D3D4B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D3D4B_din         : t_TPAR_73_DATA;
  signal TPAR_D3D4B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D3D4B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D3D4B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D3D4B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D3D4C_start                   : std_logic;
  signal TPAR_D3D4C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D3D4C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D3D4C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D3D4C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D3D4C_wea          : t_TPAR_73_1b;
  signal TPAR_D3D4C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D3D4C_din         : t_TPAR_73_DATA;
  signal TPAR_D3D4C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D3D4C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D3D4C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D3D4C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_D3D4D_start                   : std_logic;
  signal TPAR_D3D4D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_D3D4D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_D3D4D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_D3D4D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_D3D4D_wea          : t_TPAR_73_1b;
  signal TPAR_D3D4D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_D3D4D_din         : t_TPAR_73_DATA;
  signal TPAR_D3D4D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_D3D4D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_D3D4D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_D3D4D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1A_start                   : std_logic;
  signal TPAR_L1D1A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1A_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1A_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1B_start                   : std_logic;
  signal TPAR_L1D1B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1B_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1B_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1C_start                   : std_logic;
  signal TPAR_L1D1C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1C_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1C_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1D_start                   : std_logic;
  signal TPAR_L1D1D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1D_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1D_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1E_start                   : std_logic;
  signal TPAR_L1D1E_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1E_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1E_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1E_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1E_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1E_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1E_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1E_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1E_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1E_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1E_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1F_start                   : std_logic;
  signal TPAR_L1D1F_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1F_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1F_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1F_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1F_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1F_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1F_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1F_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1F_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1F_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1F_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1G_start                   : std_logic;
  signal TPAR_L1D1G_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1G_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1G_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1G_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1G_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1G_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1G_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1G_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1G_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1G_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1G_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L1D1H_start                   : std_logic;
  signal TPAR_L1D1H_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L1D1H_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L1D1H_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L1D1H_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L1D1H_wea          : t_TPAR_73_1b;
  signal TPAR_L1D1H_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L1D1H_din         : t_TPAR_73_DATA;
  signal TPAR_L1D1H_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L1D1H_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L1D1H_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L1D1H_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2D1A_start                   : std_logic;
  signal TPAR_L2D1A_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2D1A_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2D1A_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2D1A_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2D1A_wea          : t_TPAR_73_1b;
  signal TPAR_L2D1A_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2D1A_din         : t_TPAR_73_DATA;
  signal TPAR_L2D1A_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2D1A_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2D1A_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2D1A_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2D1B_start                   : std_logic;
  signal TPAR_L2D1B_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2D1B_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2D1B_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2D1B_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2D1B_wea          : t_TPAR_73_1b;
  signal TPAR_L2D1B_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2D1B_din         : t_TPAR_73_DATA;
  signal TPAR_L2D1B_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2D1B_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2D1B_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2D1B_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2D1C_start                   : std_logic;
  signal TPAR_L2D1C_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2D1C_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2D1C_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2D1C_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2D1C_wea          : t_TPAR_73_1b;
  signal TPAR_L2D1C_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2D1C_din         : t_TPAR_73_DATA;
  signal TPAR_L2D1C_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2D1C_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2D1C_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2D1C_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal TPAR_L2D1D_start                   : std_logic;
  signal TPAR_L2D1D_wea_delay          : t_TPAR_73_1b;
  signal TPAR_L2D1D_writeaddr_delay   : t_TPAR_73_ADDR;
  signal TPAR_L2D1D_din_delay         : t_TPAR_73_DATA;
  signal TPAR_L2D1D_dummy   : std_logic_vector(1 downto 0);
  signal TPAR_L2D1D_wea          : t_TPAR_73_1b;
  signal TPAR_L2D1D_writeaddr   : t_TPAR_73_ADDR;
  signal TPAR_L2D1D_din         : t_TPAR_73_DATA;
  signal TPAR_L2D1D_enb          : t_TPAR_73_1b := '1';
  --signal TPAR_L2D1D_V_readaddr    : t_TPAR_73_ADDR;
  --signal TPAR_L2D1D_V_dout        : t_TPAR_73_DATA;
  --signal TPAR_L2D1D_AV_dout_nent  : t_TPAR_73_NENT; -- (#page)
  signal IR_PS10G_1_A_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_1_A_start : std_logic := '0';
  signal IR_PS10G_1_B_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_1_B_start : std_logic := '0';
  signal IR_PS10G_2_A_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_2_A_start : std_logic := '0';
  signal IR_PS10G_2_B_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_2_B_start : std_logic := '0';
  signal IR_PS10G_3_A_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_3_A_start : std_logic := '0';
  signal IR_PS10G_3_B_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_3_B_start : std_logic := '0';
  signal IR_PS10G_4_A_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_4_A_start : std_logic := '0';
  signal IR_PS10G_4_B_bx : std_logic_vector(2 downto 0);
  signal IR_PS10G_4_B_start : std_logic := '0';
  signal IR_PS_1_A_bx : std_logic_vector(2 downto 0);
  signal IR_PS_1_A_start : std_logic := '0';
  signal IR_PS_1_B_bx : std_logic_vector(2 downto 0);
  signal IR_PS_1_B_start : std_logic := '0';
  signal IR_PS_2_A_bx : std_logic_vector(2 downto 0);
  signal IR_PS_2_A_start : std_logic := '0';
  signal IR_PS_2_B_bx : std_logic_vector(2 downto 0);
  signal IR_PS_2_B_start : std_logic := '0';
  signal IR_negPS10G_1_A_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_1_A_start : std_logic := '0';
  signal IR_negPS10G_1_B_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_1_B_start : std_logic := '0';
  signal IR_negPS10G_2_A_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_2_A_start : std_logic := '0';
  signal IR_negPS10G_2_B_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_2_B_start : std_logic := '0';
  signal IR_negPS10G_3_A_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_3_A_start : std_logic := '0';
  signal IR_negPS10G_3_B_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_3_B_start : std_logic := '0';
  signal IR_negPS10G_4_A_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_4_A_start : std_logic := '0';
  signal IR_negPS10G_4_B_bx : std_logic_vector(2 downto 0);
  signal IR_negPS10G_4_B_start : std_logic := '0';
  signal IR_negPS_1_A_bx : std_logic_vector(2 downto 0);
  signal IR_negPS_1_A_start : std_logic := '0';
  signal IR_negPS_1_B_bx : std_logic_vector(2 downto 0);
  signal IR_negPS_1_B_start : std_logic := '0';
  signal IR_negPS_2_A_bx : std_logic_vector(2 downto 0);
  signal IR_negPS_2_A_start : std_logic := '0';
  signal IR_negPS_2_B_bx : std_logic_vector(2 downto 0);
  signal IR_negPS_2_B_start : std_logic := '0';
  signal IR_2S_1_A_bx : std_logic_vector(2 downto 0);
  signal IR_2S_1_A_start : std_logic := '0';
  signal IR_2S_1_B_bx : std_logic_vector(2 downto 0);
  signal IR_2S_1_B_start : std_logic := '0';
  signal IR_2S_2_A_bx : std_logic_vector(2 downto 0);
  signal IR_2S_2_A_start : std_logic := '0';
  signal IR_2S_2_B_bx : std_logic_vector(2 downto 0);
  signal IR_2S_2_B_start : std_logic := '0';
  signal IR_2S_3_A_bx : std_logic_vector(2 downto 0);
  signal IR_2S_3_A_start : std_logic := '0';
  signal IR_2S_3_B_bx : std_logic_vector(2 downto 0);
  signal IR_2S_3_B_start : std_logic := '0';
  signal IR_2S_4_A_bx : std_logic_vector(2 downto 0);
  signal IR_2S_4_A_start : std_logic := '0';
  signal IR_2S_4_B_bx : std_logic_vector(2 downto 0);
  signal IR_2S_4_B_start : std_logic := '0';
  signal IR_2S_5_A_bx : std_logic_vector(2 downto 0);
  signal IR_2S_5_A_start : std_logic := '0';
  signal IR_2S_5_B_bx : std_logic_vector(2 downto 0);
  signal IR_2S_5_B_start : std_logic := '0';
  signal IR_2S_6_A_bx : std_logic_vector(2 downto 0);
  signal IR_2S_6_A_start : std_logic := '0';
  signal IR_2S_6_B_bx : std_logic_vector(2 downto 0);
  signal IR_2S_6_B_start : std_logic := '0';
  signal IR_neg2S_1_A_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_1_A_start : std_logic := '0';
  signal IR_neg2S_1_B_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_1_B_start : std_logic := '0';
  signal IR_neg2S_2_A_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_2_A_start : std_logic := '0';
  signal IR_neg2S_2_B_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_2_B_start : std_logic := '0';
  signal IR_neg2S_3_A_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_3_A_start : std_logic := '0';
  signal IR_neg2S_3_B_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_3_B_start : std_logic := '0';
  signal IR_neg2S_4_A_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_4_A_start : std_logic := '0';
  signal IR_neg2S_4_B_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_4_B_start : std_logic := '0';
  signal IR_neg2S_5_A_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_5_A_start : std_logic := '0';
  signal IR_neg2S_5_B_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_5_B_start : std_logic := '0';
  signal IR_neg2S_6_A_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_6_A_start : std_logic := '0';
  signal IR_neg2S_6_B_bx : std_logic_vector(2 downto 0);
  signal IR_neg2S_6_B_start : std_logic := '0';
  signal IR_done : std_logic := '0';
  signal IR_bx_out : std_logic_vector(2 downto 0);
  signal IR_bx_out_vld : std_logic;
  signal VMR_L1PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHIA_start : std_logic := '0';
  signal VMR_L1PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHIB_start : std_logic := '0';
  signal VMR_L1PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHIC_start : std_logic := '0';
  signal VMR_L1PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHID_start : std_logic := '0';
  signal VMR_L1PHIE_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHIE_start : std_logic := '0';
  signal VMR_L1PHIF_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHIF_start : std_logic := '0';
  signal VMR_L1PHIG_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHIG_start : std_logic := '0';
  signal VMR_L1PHIH_bx : std_logic_vector(2 downto 0);
  signal VMR_L1PHIH_start : std_logic := '0';
  signal VMR_L2PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_L2PHIA_start : std_logic := '0';
  signal VMR_L2PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_L2PHIB_start : std_logic := '0';
  signal VMR_L2PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_L2PHIC_start : std_logic := '0';
  signal VMR_L2PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_L2PHID_start : std_logic := '0';
  signal VMR_L3PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_L3PHIA_start : std_logic := '0';
  signal VMR_L3PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_L3PHIB_start : std_logic := '0';
  signal VMR_L3PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_L3PHIC_start : std_logic := '0';
  signal VMR_L3PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_L3PHID_start : std_logic := '0';
  signal VMR_L4PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_L4PHIA_start : std_logic := '0';
  signal VMR_L4PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_L4PHIB_start : std_logic := '0';
  signal VMR_L4PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_L4PHIC_start : std_logic := '0';
  signal VMR_L4PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_L4PHID_start : std_logic := '0';
  signal VMR_L5PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_L5PHIA_start : std_logic := '0';
  signal VMR_L5PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_L5PHIB_start : std_logic := '0';
  signal VMR_L5PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_L5PHIC_start : std_logic := '0';
  signal VMR_L5PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_L5PHID_start : std_logic := '0';
  signal VMR_L6PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_L6PHIA_start : std_logic := '0';
  signal VMR_L6PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_L6PHIB_start : std_logic := '0';
  signal VMR_L6PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_L6PHIC_start : std_logic := '0';
  signal VMR_L6PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_L6PHID_start : std_logic := '0';
  signal VMR_D1PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_D1PHIA_start : std_logic := '0';
  signal VMR_D1PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_D1PHIB_start : std_logic := '0';
  signal VMR_D1PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_D1PHIC_start : std_logic := '0';
  signal VMR_D1PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_D1PHID_start : std_logic := '0';
  signal VMR_D2PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_D2PHIA_start : std_logic := '0';
  signal VMR_D2PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_D2PHIB_start : std_logic := '0';
  signal VMR_D2PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_D2PHIC_start : std_logic := '0';
  signal VMR_D2PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_D2PHID_start : std_logic := '0';
  signal VMR_D3PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_D3PHIA_start : std_logic := '0';
  signal VMR_D3PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_D3PHIB_start : std_logic := '0';
  signal VMR_D3PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_D3PHIC_start : std_logic := '0';
  signal VMR_D3PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_D3PHID_start : std_logic := '0';
  signal VMR_D4PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_D4PHIA_start : std_logic := '0';
  signal VMR_D4PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_D4PHIB_start : std_logic := '0';
  signal VMR_D4PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_D4PHIC_start : std_logic := '0';
  signal VMR_D4PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_D4PHID_start : std_logic := '0';
  signal VMR_D5PHIA_bx : std_logic_vector(2 downto 0);
  signal VMR_D5PHIA_start : std_logic := '0';
  signal VMR_D5PHIB_bx : std_logic_vector(2 downto 0);
  signal VMR_D5PHIB_start : std_logic := '0';
  signal VMR_D5PHIC_bx : std_logic_vector(2 downto 0);
  signal VMR_D5PHIC_start : std_logic := '0';
  signal VMR_D5PHID_bx : std_logic_vector(2 downto 0);
  signal VMR_D5PHID_start : std_logic := '0';
  signal VMR_done : std_logic := '0';
  signal VMR_bx_out : std_logic_vector(2 downto 0);
  signal VMR_bx_out_vld : std_logic;
  signal TP_L1L2A_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2A_start : std_logic := '0';
  signal TP_L1L2B_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2B_start : std_logic := '0';
  signal TP_L1L2C_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2C_start : std_logic := '0';
  signal TP_L1L2D_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2D_start : std_logic := '0';
  signal TP_L1L2E_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2E_start : std_logic := '0';
  signal TP_L1L2F_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2F_start : std_logic := '0';
  signal TP_L1L2G_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2G_start : std_logic := '0';
  signal TP_L1L2H_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2H_start : std_logic := '0';
  signal TP_L1L2I_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2I_start : std_logic := '0';
  signal TP_L1L2J_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2J_start : std_logic := '0';
  signal TP_L1L2K_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2K_start : std_logic := '0';
  signal TP_L1L2L_bx : std_logic_vector(2 downto 0);
  signal TP_L1L2L_start : std_logic := '0';
  signal TP_L2L3A_bx : std_logic_vector(2 downto 0);
  signal TP_L2L3A_start : std_logic := '0';
  signal TP_L2L3B_bx : std_logic_vector(2 downto 0);
  signal TP_L2L3B_start : std_logic := '0';
  signal TP_L2L3C_bx : std_logic_vector(2 downto 0);
  signal TP_L2L3C_start : std_logic := '0';
  signal TP_L2L3D_bx : std_logic_vector(2 downto 0);
  signal TP_L2L3D_start : std_logic := '0';
  signal TP_L3L4A_bx : std_logic_vector(2 downto 0);
  signal TP_L3L4A_start : std_logic := '0';
  signal TP_L3L4B_bx : std_logic_vector(2 downto 0);
  signal TP_L3L4B_start : std_logic := '0';
  signal TP_L3L4C_bx : std_logic_vector(2 downto 0);
  signal TP_L3L4C_start : std_logic := '0';
  signal TP_L3L4D_bx : std_logic_vector(2 downto 0);
  signal TP_L3L4D_start : std_logic := '0';
  signal TP_L5L6A_bx : std_logic_vector(2 downto 0);
  signal TP_L5L6A_start : std_logic := '0';
  signal TP_L5L6B_bx : std_logic_vector(2 downto 0);
  signal TP_L5L6B_start : std_logic := '0';
  signal TP_L5L6C_bx : std_logic_vector(2 downto 0);
  signal TP_L5L6C_start : std_logic := '0';
  signal TP_L5L6D_bx : std_logic_vector(2 downto 0);
  signal TP_L5L6D_start : std_logic := '0';
  signal TP_D1D2A_bx : std_logic_vector(2 downto 0);
  signal TP_D1D2A_start : std_logic := '0';
  signal TP_D1D2B_bx : std_logic_vector(2 downto 0);
  signal TP_D1D2B_start : std_logic := '0';
  signal TP_D1D2C_bx : std_logic_vector(2 downto 0);
  signal TP_D1D2C_start : std_logic := '0';
  signal TP_D1D2D_bx : std_logic_vector(2 downto 0);
  signal TP_D1D2D_start : std_logic := '0';
  signal TP_D3D4A_bx : std_logic_vector(2 downto 0);
  signal TP_D3D4A_start : std_logic := '0';
  signal TP_D3D4B_bx : std_logic_vector(2 downto 0);
  signal TP_D3D4B_start : std_logic := '0';
  signal TP_D3D4C_bx : std_logic_vector(2 downto 0);
  signal TP_D3D4C_start : std_logic := '0';
  signal TP_D3D4D_bx : std_logic_vector(2 downto 0);
  signal TP_D3D4D_start : std_logic := '0';
  signal TP_L1D1A_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1A_start : std_logic := '0';
  signal TP_L1D1B_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1B_start : std_logic := '0';
  signal TP_L1D1C_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1C_start : std_logic := '0';
  signal TP_L1D1D_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1D_start : std_logic := '0';
  signal TP_L1D1E_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1E_start : std_logic := '0';
  signal TP_L1D1F_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1F_start : std_logic := '0';
  signal TP_L1D1G_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1G_start : std_logic := '0';
  signal TP_L1D1H_bx : std_logic_vector(2 downto 0);
  signal TP_L1D1H_start : std_logic := '0';
  signal TP_L2D1A_bx : std_logic_vector(2 downto 0);
  signal TP_L2D1A_start : std_logic := '0';
  signal TP_L2D1B_bx : std_logic_vector(2 downto 0);
  signal TP_L2D1B_start : std_logic := '0';
  signal TP_L2D1C_bx : std_logic_vector(2 downto 0);
  signal TP_L2D1C_start : std_logic := '0';
  signal TP_L2D1D_bx : std_logic_vector(2 downto 0);
  signal TP_L2D1D_start : std_logic := '0';

  --signal AS_D1PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D1PHIAn1_bx_vld : std_logic;
  --signal AS_D1PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D1PHIBn1_bx_vld : std_logic;
  --signal AS_D1PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D1PHICn1_bx_vld : std_logic;
  --signal AS_D1PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D1PHIDn1_bx_vld : std_logic;
  --signal AS_D2PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D2PHIAn1_bx_vld : std_logic;
  --signal AS_D2PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D2PHIBn1_bx_vld : std_logic;
  --signal AS_D2PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D2PHICn1_bx_vld : std_logic;
  --signal AS_D2PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D2PHIDn1_bx_vld : std_logic;
  --signal AS_D3PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D3PHIAn1_bx_vld : std_logic;
  --signal AS_D3PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D3PHIBn1_bx_vld : std_logic;
  --signal AS_D3PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D3PHICn1_bx_vld : std_logic;
  --signal AS_D3PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D3PHIDn1_bx_vld : std_logic;
  --signal AS_D4PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D4PHIAn1_bx_vld : std_logic;
  --signal AS_D4PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D4PHIBn1_bx_vld : std_logic;
  --signal AS_D4PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D4PHICn1_bx_vld : std_logic;
  --signal AS_D4PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D4PHIDn1_bx_vld : std_logic;
  --signal AS_D5PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D5PHIAn1_bx_vld : std_logic;
  --signal AS_D5PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D5PHIBn1_bx_vld : std_logic;
  --signal AS_D5PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D5PHICn1_bx_vld : std_logic;
  --signal AS_D5PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_D5PHIDn1_bx_vld : std_logic;
  --signal AS_L1PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHIAn1_bx_vld : std_logic;
  --signal AS_L1PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHIBn1_bx_vld : std_logic;
  --signal AS_L1PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHICn1_bx_vld : std_logic;
  --signal AS_L1PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHIDn1_bx_vld : std_logic;
  --signal AS_L1PHIEn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHIEn1_bx_vld : std_logic;
  --signal AS_L1PHIFn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHIFn1_bx_vld : std_logic;
  --signal AS_L1PHIGn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHIGn1_bx_vld : std_logic;
  --signal AS_L1PHIHn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L1PHIHn1_bx_vld : std_logic;
  --signal AS_L2PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L2PHIAn1_bx_vld : std_logic;
  --signal AS_L2PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L2PHIBn1_bx_vld : std_logic;
  --signal AS_L2PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L2PHICn1_bx_vld : std_logic;
  --signal AS_L2PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L2PHIDn1_bx_vld : std_logic;
  --signal AS_L3PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L3PHIAn1_bx_vld : std_logic;
  --signal AS_L3PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L3PHIBn1_bx_vld : std_logic;
  --signal AS_L3PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L3PHICn1_bx_vld : std_logic;
  --signal AS_L3PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L3PHIDn1_bx_vld : std_logic;
  --signal AS_L4PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L4PHIAn1_bx_vld : std_logic;
  --signal AS_L4PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L4PHIBn1_bx_vld : std_logic;
  --signal AS_L4PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L4PHICn1_bx_vld : std_logic;
  --signal AS_L4PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L4PHIDn1_bx_vld : std_logic;
  --signal AS_L5PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L5PHIAn1_bx_vld : std_logic;
  --signal AS_L5PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L5PHIBn1_bx_vld : std_logic;
  --signal AS_L5PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L5PHICn1_bx_vld : std_logic;
  --signal AS_L5PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L5PHIDn1_bx_vld : std_logic;
  --signal AS_L6PHIAn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L6PHIAn1_bx_vld : std_logic;
  --signal AS_L6PHIBn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L6PHIBn1_bx_vld : std_logic;
  --signal AS_L6PHICn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L6PHICn1_bx_vld : std_logic;
  --signal AS_L6PHIDn1_bx : std_logic_vector(2 downto 0);
  --signal AS_L6PHIDn1_bx_vld : std_logic;
  --signal TPARD1D2ABCD_bx : std_logic_vector(2 downto 0);
  --signal TPARD1D2ABCD_bx_vld : std_logic;
  --signal TPARD3D4ABCD_bx : std_logic_vector(2 downto 0);
  --signal TPARD3D4ABCD_bx_vld : std_logic;
  --signal TPARL1D1ABCD_bx : std_logic_vector(2 downto 0);
  --signal TPARL1D1ABCD_bx_vld : std_logic;
  --signal TPARL1D1EFGH_bx : std_logic_vector(2 downto 0);
  --signal TPARL1D1EFGH_bx_vld : std_logic;
  --signal TPARL1L2ABC_bx : std_logic_vector(2 downto 0);
  --signal TPARL1L2ABC_bx_vld : std_logic;
  --signal TPARL1L2DE_bx : std_logic_vector(2 downto 0);
  --signal TPARL1L2DE_bx_vld : std_logic;
  --signal TPARL1L2F_bx : std_logic_vector(2 downto 0);
  --signal TPARL1L2F_bx_vld : std_logic;
  --signal TPARL1L2G_bx : std_logic_vector(2 downto 0);
  --signal TPARL1L2G_bx_vld : std_logic;
  --signal TPARL1L2HI_bx : std_logic_vector(2 downto 0);
  --signal TPARL1L2HI_bx_vld : std_logic;
  --signal TPARL1L2JKL_bx : std_logic_vector(2 downto 0);
  --signal TPARL1L2JKL_bx_vld : std_logic;
  --signal TPARL2D1ABCD_bx : std_logic_vector(2 downto 0);
  --signal TPARL2D1ABCD_bx_vld : std_logic;
  --signal TPARL2L3ABCD_bx : std_logic_vector(2 downto 0);
  --signal TPARL2L3ABCD_bx_vld : std_logic;
  --signal TPARL3L4AB_bx : std_logic_vector(2 downto 0);
  --signal TPARL3L4AB_bx_vld : std_logic;
  --signal TPARL3L4CD_bx : std_logic_vector(2 downto 0);
  --signal TPARL3L4CD_bx_vld : std_logic;
  --signal TPARL5L6ABCD_bx : std_logic_vector(2 downto 0);
  --signal TPARL5L6ABCD_bx_vld : std_logic;

begin

    IL_L1PHIA_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIA_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIA_PS10G_1_A_wea_delay,
        addra     => IL_L1PHIA_PS10G_1_A_writeaddr_delay,
        dina      => IL_L1PHIA_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIA_PS10G_1_A_V_readaddr,
        doutb     => IL_L1PHIA_PS10G_1_A_V_dout,
        sync_nent => IL_L1PHIA_PS10G_1_A_start,
        nent_o    => IL_L1PHIA_PS10G_1_A_AV_dout_nent
      );

    IL_L1PHIA_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIA_PS10G_1_A_wea,
        addra     => IL_L1PHIA_PS10G_1_A_writeaddr,
        dina      => IL_L1PHIA_PS10G_1_A_din,
        wea_out       => IL_L1PHIA_PS10G_1_A_wea_delay,
        addra_out     => IL_L1PHIA_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_L1PHIA_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIA_PS10G_1_A_start
      );

    IL_L1PHIB_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIB_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIB_PS10G_1_A_wea_delay,
        addra     => IL_L1PHIB_PS10G_1_A_writeaddr_delay,
        dina      => IL_L1PHIB_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIB_PS10G_1_A_V_readaddr,
        doutb     => IL_L1PHIB_PS10G_1_A_V_dout,
        sync_nent => IL_L1PHIB_PS10G_1_A_start,
        nent_o    => IL_L1PHIB_PS10G_1_A_AV_dout_nent
      );

    IL_L1PHIB_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIB_PS10G_1_A_wea,
        addra     => IL_L1PHIB_PS10G_1_A_writeaddr,
        dina      => IL_L1PHIB_PS10G_1_A_din,
        wea_out       => IL_L1PHIB_PS10G_1_A_wea_delay,
        addra_out     => IL_L1PHIB_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_L1PHIB_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIB_PS10G_1_A_start
      );

    IL_L1PHIC_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIC_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIC_PS10G_1_A_wea_delay,
        addra     => IL_L1PHIC_PS10G_1_A_writeaddr_delay,
        dina      => IL_L1PHIC_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIC_PS10G_1_A_V_readaddr,
        doutb     => IL_L1PHIC_PS10G_1_A_V_dout,
        sync_nent => IL_L1PHIC_PS10G_1_A_start,
        nent_o    => IL_L1PHIC_PS10G_1_A_AV_dout_nent
      );

    IL_L1PHIC_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIC_PS10G_1_A_wea,
        addra     => IL_L1PHIC_PS10G_1_A_writeaddr,
        dina      => IL_L1PHIC_PS10G_1_A_din,
        wea_out       => IL_L1PHIC_PS10G_1_A_wea_delay,
        addra_out     => IL_L1PHIC_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_L1PHIC_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIC_PS10G_1_A_start
      );

    IL_L1PHID_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHID_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHID_PS10G_1_A_wea_delay,
        addra     => IL_L1PHID_PS10G_1_A_writeaddr_delay,
        dina      => IL_L1PHID_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHID_PS10G_1_A_V_readaddr,
        doutb     => IL_L1PHID_PS10G_1_A_V_dout,
        sync_nent => IL_L1PHID_PS10G_1_A_start,
        nent_o    => IL_L1PHID_PS10G_1_A_AV_dout_nent
      );

    IL_L1PHID_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHID_PS10G_1_A_wea,
        addra     => IL_L1PHID_PS10G_1_A_writeaddr,
        dina      => IL_L1PHID_PS10G_1_A_din,
        wea_out       => IL_L1PHID_PS10G_1_A_wea_delay,
        addra_out     => IL_L1PHID_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_L1PHID_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHID_PS10G_1_A_start
      );

    IL_L1PHIE_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIE_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIE_PS10G_1_A_wea_delay,
        addra     => IL_L1PHIE_PS10G_1_A_writeaddr_delay,
        dina      => IL_L1PHIE_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIE_PS10G_1_A_V_readaddr,
        doutb     => IL_L1PHIE_PS10G_1_A_V_dout,
        sync_nent => IL_L1PHIE_PS10G_1_A_start,
        nent_o    => IL_L1PHIE_PS10G_1_A_AV_dout_nent
      );

    IL_L1PHIE_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIE_PS10G_1_A_wea,
        addra     => IL_L1PHIE_PS10G_1_A_writeaddr,
        dina      => IL_L1PHIE_PS10G_1_A_din,
        wea_out       => IL_L1PHIE_PS10G_1_A_wea_delay,
        addra_out     => IL_L1PHIE_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_L1PHIE_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIE_PS10G_1_A_start
      );

    IL_L1PHIG_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIG_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIG_PS10G_1_B_wea_delay,
        addra     => IL_L1PHIG_PS10G_1_B_writeaddr_delay,
        dina      => IL_L1PHIG_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIG_PS10G_1_B_V_readaddr,
        doutb     => IL_L1PHIG_PS10G_1_B_V_dout,
        sync_nent => IL_L1PHIG_PS10G_1_B_start,
        nent_o    => IL_L1PHIG_PS10G_1_B_AV_dout_nent
      );

    IL_L1PHIG_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIG_PS10G_1_B_wea,
        addra     => IL_L1PHIG_PS10G_1_B_writeaddr,
        dina      => IL_L1PHIG_PS10G_1_B_din,
        wea_out       => IL_L1PHIG_PS10G_1_B_wea_delay,
        addra_out     => IL_L1PHIG_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_L1PHIG_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIG_PS10G_1_B_start
      );

    IL_L1PHIH_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIH_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIH_PS10G_1_B_wea_delay,
        addra     => IL_L1PHIH_PS10G_1_B_writeaddr_delay,
        dina      => IL_L1PHIH_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIH_PS10G_1_B_V_readaddr,
        doutb     => IL_L1PHIH_PS10G_1_B_V_dout,
        sync_nent => IL_L1PHIH_PS10G_1_B_start,
        nent_o    => IL_L1PHIH_PS10G_1_B_AV_dout_nent
      );

    IL_L1PHIH_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIH_PS10G_1_B_wea,
        addra     => IL_L1PHIH_PS10G_1_B_writeaddr,
        dina      => IL_L1PHIH_PS10G_1_B_din,
        wea_out       => IL_L1PHIH_PS10G_1_B_wea_delay,
        addra_out     => IL_L1PHIH_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_L1PHIH_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIH_PS10G_1_B_start
      );

    IL_D1PHIA_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIA_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIA_PS10G_1_A_wea_delay,
        addra     => IL_D1PHIA_PS10G_1_A_writeaddr_delay,
        dina      => IL_D1PHIA_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIA_PS10G_1_A_V_readaddr,
        doutb     => IL_D1PHIA_PS10G_1_A_V_dout,
        sync_nent => IL_D1PHIA_PS10G_1_A_start,
        nent_o    => IL_D1PHIA_PS10G_1_A_AV_dout_nent
      );

    IL_D1PHIA_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIA_PS10G_1_A_wea,
        addra     => IL_D1PHIA_PS10G_1_A_writeaddr,
        dina      => IL_D1PHIA_PS10G_1_A_din,
        wea_out       => IL_D1PHIA_PS10G_1_A_wea_delay,
        addra_out     => IL_D1PHIA_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D1PHIA_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIA_PS10G_1_A_start
      );

    IL_D1PHIB_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_PS10G_1_A_wea_delay,
        addra     => IL_D1PHIB_PS10G_1_A_writeaddr_delay,
        dina      => IL_D1PHIB_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_PS10G_1_A_V_readaddr,
        doutb     => IL_D1PHIB_PS10G_1_A_V_dout,
        sync_nent => IL_D1PHIB_PS10G_1_A_start,
        nent_o    => IL_D1PHIB_PS10G_1_A_AV_dout_nent
      );

    IL_D1PHIB_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_PS10G_1_A_wea,
        addra     => IL_D1PHIB_PS10G_1_A_writeaddr,
        dina      => IL_D1PHIB_PS10G_1_A_din,
        wea_out       => IL_D1PHIB_PS10G_1_A_wea_delay,
        addra_out     => IL_D1PHIB_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D1PHIB_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_PS10G_1_A_start
      );

    IL_D1PHIB_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_PS10G_1_B_wea_delay,
        addra     => IL_D1PHIB_PS10G_1_B_writeaddr_delay,
        dina      => IL_D1PHIB_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_PS10G_1_B_V_readaddr,
        doutb     => IL_D1PHIB_PS10G_1_B_V_dout,
        sync_nent => IL_D1PHIB_PS10G_1_B_start,
        nent_o    => IL_D1PHIB_PS10G_1_B_AV_dout_nent
      );

    IL_D1PHIB_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_PS10G_1_B_wea,
        addra     => IL_D1PHIB_PS10G_1_B_writeaddr,
        dina      => IL_D1PHIB_PS10G_1_B_din,
        wea_out       => IL_D1PHIB_PS10G_1_B_wea_delay,
        addra_out     => IL_D1PHIB_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D1PHIB_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_PS10G_1_B_start
      );

    IL_D1PHIC_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_PS10G_1_A_wea_delay,
        addra     => IL_D1PHIC_PS10G_1_A_writeaddr_delay,
        dina      => IL_D1PHIC_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_PS10G_1_A_V_readaddr,
        doutb     => IL_D1PHIC_PS10G_1_A_V_dout,
        sync_nent => IL_D1PHIC_PS10G_1_A_start,
        nent_o    => IL_D1PHIC_PS10G_1_A_AV_dout_nent
      );

    IL_D1PHIC_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_PS10G_1_A_wea,
        addra     => IL_D1PHIC_PS10G_1_A_writeaddr,
        dina      => IL_D1PHIC_PS10G_1_A_din,
        wea_out       => IL_D1PHIC_PS10G_1_A_wea_delay,
        addra_out     => IL_D1PHIC_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D1PHIC_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_PS10G_1_A_start
      );

    IL_D1PHIC_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_PS10G_1_B_wea_delay,
        addra     => IL_D1PHIC_PS10G_1_B_writeaddr_delay,
        dina      => IL_D1PHIC_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_PS10G_1_B_V_readaddr,
        doutb     => IL_D1PHIC_PS10G_1_B_V_dout,
        sync_nent => IL_D1PHIC_PS10G_1_B_start,
        nent_o    => IL_D1PHIC_PS10G_1_B_AV_dout_nent
      );

    IL_D1PHIC_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_PS10G_1_B_wea,
        addra     => IL_D1PHIC_PS10G_1_B_writeaddr,
        dina      => IL_D1PHIC_PS10G_1_B_din,
        wea_out       => IL_D1PHIC_PS10G_1_B_wea_delay,
        addra_out     => IL_D1PHIC_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D1PHIC_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_PS10G_1_B_start
      );

    IL_D1PHID_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHID_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHID_PS10G_1_B_wea_delay,
        addra     => IL_D1PHID_PS10G_1_B_writeaddr_delay,
        dina      => IL_D1PHID_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHID_PS10G_1_B_V_readaddr,
        doutb     => IL_D1PHID_PS10G_1_B_V_dout,
        sync_nent => IL_D1PHID_PS10G_1_B_start,
        nent_o    => IL_D1PHID_PS10G_1_B_AV_dout_nent
      );

    IL_D1PHID_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHID_PS10G_1_B_wea,
        addra     => IL_D1PHID_PS10G_1_B_writeaddr,
        dina      => IL_D1PHID_PS10G_1_B_din,
        wea_out       => IL_D1PHID_PS10G_1_B_wea_delay,
        addra_out     => IL_D1PHID_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D1PHID_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHID_PS10G_1_B_start
      );

    IL_D3PHIA_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIA_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIA_PS10G_1_A_wea_delay,
        addra     => IL_D3PHIA_PS10G_1_A_writeaddr_delay,
        dina      => IL_D3PHIA_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIA_PS10G_1_A_V_readaddr,
        doutb     => IL_D3PHIA_PS10G_1_A_V_dout,
        sync_nent => IL_D3PHIA_PS10G_1_A_start,
        nent_o    => IL_D3PHIA_PS10G_1_A_AV_dout_nent
      );

    IL_D3PHIA_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIA_PS10G_1_A_wea,
        addra     => IL_D3PHIA_PS10G_1_A_writeaddr,
        dina      => IL_D3PHIA_PS10G_1_A_din,
        wea_out       => IL_D3PHIA_PS10G_1_A_wea_delay,
        addra_out     => IL_D3PHIA_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D3PHIA_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIA_PS10G_1_A_start
      );

    IL_D3PHIB_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_PS10G_1_A_wea_delay,
        addra     => IL_D3PHIB_PS10G_1_A_writeaddr_delay,
        dina      => IL_D3PHIB_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_PS10G_1_A_V_readaddr,
        doutb     => IL_D3PHIB_PS10G_1_A_V_dout,
        sync_nent => IL_D3PHIB_PS10G_1_A_start,
        nent_o    => IL_D3PHIB_PS10G_1_A_AV_dout_nent
      );

    IL_D3PHIB_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_PS10G_1_A_wea,
        addra     => IL_D3PHIB_PS10G_1_A_writeaddr,
        dina      => IL_D3PHIB_PS10G_1_A_din,
        wea_out       => IL_D3PHIB_PS10G_1_A_wea_delay,
        addra_out     => IL_D3PHIB_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D3PHIB_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_PS10G_1_A_start
      );

    IL_D3PHIB_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_PS10G_1_B_wea_delay,
        addra     => IL_D3PHIB_PS10G_1_B_writeaddr_delay,
        dina      => IL_D3PHIB_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_PS10G_1_B_V_readaddr,
        doutb     => IL_D3PHIB_PS10G_1_B_V_dout,
        sync_nent => IL_D3PHIB_PS10G_1_B_start,
        nent_o    => IL_D3PHIB_PS10G_1_B_AV_dout_nent
      );

    IL_D3PHIB_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_PS10G_1_B_wea,
        addra     => IL_D3PHIB_PS10G_1_B_writeaddr,
        dina      => IL_D3PHIB_PS10G_1_B_din,
        wea_out       => IL_D3PHIB_PS10G_1_B_wea_delay,
        addra_out     => IL_D3PHIB_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D3PHIB_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_PS10G_1_B_start
      );

    IL_D3PHIC_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_PS10G_1_A_wea_delay,
        addra     => IL_D3PHIC_PS10G_1_A_writeaddr_delay,
        dina      => IL_D3PHIC_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_PS10G_1_A_V_readaddr,
        doutb     => IL_D3PHIC_PS10G_1_A_V_dout,
        sync_nent => IL_D3PHIC_PS10G_1_A_start,
        nent_o    => IL_D3PHIC_PS10G_1_A_AV_dout_nent
      );

    IL_D3PHIC_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_PS10G_1_A_wea,
        addra     => IL_D3PHIC_PS10G_1_A_writeaddr,
        dina      => IL_D3PHIC_PS10G_1_A_din,
        wea_out       => IL_D3PHIC_PS10G_1_A_wea_delay,
        addra_out     => IL_D3PHIC_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D3PHIC_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_PS10G_1_A_start
      );

    IL_D3PHIC_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_PS10G_1_B_wea_delay,
        addra     => IL_D3PHIC_PS10G_1_B_writeaddr_delay,
        dina      => IL_D3PHIC_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_PS10G_1_B_V_readaddr,
        doutb     => IL_D3PHIC_PS10G_1_B_V_dout,
        sync_nent => IL_D3PHIC_PS10G_1_B_start,
        nent_o    => IL_D3PHIC_PS10G_1_B_AV_dout_nent
      );

    IL_D3PHIC_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_PS10G_1_B_wea,
        addra     => IL_D3PHIC_PS10G_1_B_writeaddr,
        dina      => IL_D3PHIC_PS10G_1_B_din,
        wea_out       => IL_D3PHIC_PS10G_1_B_wea_delay,
        addra_out     => IL_D3PHIC_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D3PHIC_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_PS10G_1_B_start
      );

    IL_D3PHID_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHID_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHID_PS10G_1_B_wea_delay,
        addra     => IL_D3PHID_PS10G_1_B_writeaddr_delay,
        dina      => IL_D3PHID_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHID_PS10G_1_B_V_readaddr,
        doutb     => IL_D3PHID_PS10G_1_B_V_dout,
        sync_nent => IL_D3PHID_PS10G_1_B_start,
        nent_o    => IL_D3PHID_PS10G_1_B_AV_dout_nent
      );

    IL_D3PHID_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHID_PS10G_1_B_wea,
        addra     => IL_D3PHID_PS10G_1_B_writeaddr,
        dina      => IL_D3PHID_PS10G_1_B_din,
        wea_out       => IL_D3PHID_PS10G_1_B_wea_delay,
        addra_out     => IL_D3PHID_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D3PHID_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHID_PS10G_1_B_start
      );

    IL_D5PHIA_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIA_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIA_PS10G_1_A_wea_delay,
        addra     => IL_D5PHIA_PS10G_1_A_writeaddr_delay,
        dina      => IL_D5PHIA_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIA_PS10G_1_A_V_readaddr,
        doutb     => IL_D5PHIA_PS10G_1_A_V_dout,
        sync_nent => IL_D5PHIA_PS10G_1_A_start,
        nent_o    => IL_D5PHIA_PS10G_1_A_AV_dout_nent
      );

    IL_D5PHIA_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIA_PS10G_1_A_wea,
        addra     => IL_D5PHIA_PS10G_1_A_writeaddr,
        dina      => IL_D5PHIA_PS10G_1_A_din,
        wea_out       => IL_D5PHIA_PS10G_1_A_wea_delay,
        addra_out     => IL_D5PHIA_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D5PHIA_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIA_PS10G_1_A_start
      );

    IL_D5PHIB_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_PS10G_1_A_wea_delay,
        addra     => IL_D5PHIB_PS10G_1_A_writeaddr_delay,
        dina      => IL_D5PHIB_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_PS10G_1_A_V_readaddr,
        doutb     => IL_D5PHIB_PS10G_1_A_V_dout,
        sync_nent => IL_D5PHIB_PS10G_1_A_start,
        nent_o    => IL_D5PHIB_PS10G_1_A_AV_dout_nent
      );

    IL_D5PHIB_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_PS10G_1_A_wea,
        addra     => IL_D5PHIB_PS10G_1_A_writeaddr,
        dina      => IL_D5PHIB_PS10G_1_A_din,
        wea_out       => IL_D5PHIB_PS10G_1_A_wea_delay,
        addra_out     => IL_D5PHIB_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D5PHIB_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_PS10G_1_A_start
      );

    IL_D5PHIB_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_PS10G_1_B_wea_delay,
        addra     => IL_D5PHIB_PS10G_1_B_writeaddr_delay,
        dina      => IL_D5PHIB_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_PS10G_1_B_V_readaddr,
        doutb     => IL_D5PHIB_PS10G_1_B_V_dout,
        sync_nent => IL_D5PHIB_PS10G_1_B_start,
        nent_o    => IL_D5PHIB_PS10G_1_B_AV_dout_nent
      );

    IL_D5PHIB_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_PS10G_1_B_wea,
        addra     => IL_D5PHIB_PS10G_1_B_writeaddr,
        dina      => IL_D5PHIB_PS10G_1_B_din,
        wea_out       => IL_D5PHIB_PS10G_1_B_wea_delay,
        addra_out     => IL_D5PHIB_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D5PHIB_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_PS10G_1_B_start
      );

    IL_D5PHIC_PS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_PS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_PS10G_1_A_wea_delay,
        addra     => IL_D5PHIC_PS10G_1_A_writeaddr_delay,
        dina      => IL_D5PHIC_PS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_PS10G_1_A_V_readaddr,
        doutb     => IL_D5PHIC_PS10G_1_A_V_dout,
        sync_nent => IL_D5PHIC_PS10G_1_A_start,
        nent_o    => IL_D5PHIC_PS10G_1_A_AV_dout_nent
      );

    IL_D5PHIC_PS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_PS10G_1_A_wea,
        addra     => IL_D5PHIC_PS10G_1_A_writeaddr,
        dina      => IL_D5PHIC_PS10G_1_A_din,
        wea_out       => IL_D5PHIC_PS10G_1_A_wea_delay,
        addra_out     => IL_D5PHIC_PS10G_1_A_writeaddr_delay,
        dina_out      => IL_D5PHIC_PS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_PS10G_1_A_start
      );

    IL_D5PHIC_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_PS10G_1_B_wea_delay,
        addra     => IL_D5PHIC_PS10G_1_B_writeaddr_delay,
        dina      => IL_D5PHIC_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_PS10G_1_B_V_readaddr,
        doutb     => IL_D5PHIC_PS10G_1_B_V_dout,
        sync_nent => IL_D5PHIC_PS10G_1_B_start,
        nent_o    => IL_D5PHIC_PS10G_1_B_AV_dout_nent
      );

    IL_D5PHIC_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_PS10G_1_B_wea,
        addra     => IL_D5PHIC_PS10G_1_B_writeaddr,
        dina      => IL_D5PHIC_PS10G_1_B_din,
        wea_out       => IL_D5PHIC_PS10G_1_B_wea_delay,
        addra_out     => IL_D5PHIC_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D5PHIC_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_PS10G_1_B_start
      );

    IL_D5PHID_PS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHID_PS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHID_PS10G_1_B_wea_delay,
        addra     => IL_D5PHID_PS10G_1_B_writeaddr_delay,
        dina      => IL_D5PHID_PS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHID_PS10G_1_B_V_readaddr,
        doutb     => IL_D5PHID_PS10G_1_B_V_dout,
        sync_nent => IL_D5PHID_PS10G_1_B_start,
        nent_o    => IL_D5PHID_PS10G_1_B_AV_dout_nent
      );

    IL_D5PHID_PS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHID_PS10G_1_B_wea,
        addra     => IL_D5PHID_PS10G_1_B_writeaddr,
        dina      => IL_D5PHID_PS10G_1_B_din,
        wea_out       => IL_D5PHID_PS10G_1_B_wea_delay,
        addra_out     => IL_D5PHID_PS10G_1_B_writeaddr_delay,
        dina_out      => IL_D5PHID_PS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHID_PS10G_1_B_start
      );

    IL_L1PHIA_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIA_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIA_PS10G_2_A_wea_delay,
        addra     => IL_L1PHIA_PS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIA_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIA_PS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIA_PS10G_2_A_V_dout,
        sync_nent => IL_L1PHIA_PS10G_2_A_start,
        nent_o    => IL_L1PHIA_PS10G_2_A_AV_dout_nent
      );

    IL_L1PHIA_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIA_PS10G_2_A_wea,
        addra     => IL_L1PHIA_PS10G_2_A_writeaddr,
        dina      => IL_L1PHIA_PS10G_2_A_din,
        wea_out       => IL_L1PHIA_PS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIA_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIA_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIA_PS10G_2_A_start
      );

    IL_L1PHIB_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIB_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIB_PS10G_2_A_wea_delay,
        addra     => IL_L1PHIB_PS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIB_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIB_PS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIB_PS10G_2_A_V_dout,
        sync_nent => IL_L1PHIB_PS10G_2_A_start,
        nent_o    => IL_L1PHIB_PS10G_2_A_AV_dout_nent
      );

    IL_L1PHIB_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIB_PS10G_2_A_wea,
        addra     => IL_L1PHIB_PS10G_2_A_writeaddr,
        dina      => IL_L1PHIB_PS10G_2_A_din,
        wea_out       => IL_L1PHIB_PS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIB_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIB_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIB_PS10G_2_A_start
      );

    IL_L1PHIC_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIC_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIC_PS10G_2_A_wea_delay,
        addra     => IL_L1PHIC_PS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIC_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIC_PS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIC_PS10G_2_A_V_dout,
        sync_nent => IL_L1PHIC_PS10G_2_A_start,
        nent_o    => IL_L1PHIC_PS10G_2_A_AV_dout_nent
      );

    IL_L1PHIC_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIC_PS10G_2_A_wea,
        addra     => IL_L1PHIC_PS10G_2_A_writeaddr,
        dina      => IL_L1PHIC_PS10G_2_A_din,
        wea_out       => IL_L1PHIC_PS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIC_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIC_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIC_PS10G_2_A_start
      );

    IL_L1PHID_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHID_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHID_PS10G_2_A_wea_delay,
        addra     => IL_L1PHID_PS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHID_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHID_PS10G_2_A_V_readaddr,
        doutb     => IL_L1PHID_PS10G_2_A_V_dout,
        sync_nent => IL_L1PHID_PS10G_2_A_start,
        nent_o    => IL_L1PHID_PS10G_2_A_AV_dout_nent
      );

    IL_L1PHID_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHID_PS10G_2_A_wea,
        addra     => IL_L1PHID_PS10G_2_A_writeaddr,
        dina      => IL_L1PHID_PS10G_2_A_din,
        wea_out       => IL_L1PHID_PS10G_2_A_wea_delay,
        addra_out     => IL_L1PHID_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHID_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHID_PS10G_2_A_start
      );

    IL_L1PHID_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHID_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHID_PS10G_2_B_wea_delay,
        addra     => IL_L1PHID_PS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHID_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHID_PS10G_2_B_V_readaddr,
        doutb     => IL_L1PHID_PS10G_2_B_V_dout,
        sync_nent => IL_L1PHID_PS10G_2_B_start,
        nent_o    => IL_L1PHID_PS10G_2_B_AV_dout_nent
      );

    IL_L1PHID_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHID_PS10G_2_B_wea,
        addra     => IL_L1PHID_PS10G_2_B_writeaddr,
        dina      => IL_L1PHID_PS10G_2_B_din,
        wea_out       => IL_L1PHID_PS10G_2_B_wea_delay,
        addra_out     => IL_L1PHID_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHID_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHID_PS10G_2_B_start
      );

    IL_L1PHIE_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIE_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIE_PS10G_2_A_wea_delay,
        addra     => IL_L1PHIE_PS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIE_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIE_PS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIE_PS10G_2_A_V_dout,
        sync_nent => IL_L1PHIE_PS10G_2_A_start,
        nent_o    => IL_L1PHIE_PS10G_2_A_AV_dout_nent
      );

    IL_L1PHIE_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIE_PS10G_2_A_wea,
        addra     => IL_L1PHIE_PS10G_2_A_writeaddr,
        dina      => IL_L1PHIE_PS10G_2_A_din,
        wea_out       => IL_L1PHIE_PS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIE_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIE_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIE_PS10G_2_A_start
      );

    IL_L1PHIE_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIE_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIE_PS10G_2_B_wea_delay,
        addra     => IL_L1PHIE_PS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIE_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIE_PS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIE_PS10G_2_B_V_dout,
        sync_nent => IL_L1PHIE_PS10G_2_B_start,
        nent_o    => IL_L1PHIE_PS10G_2_B_AV_dout_nent
      );

    IL_L1PHIE_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIE_PS10G_2_B_wea,
        addra     => IL_L1PHIE_PS10G_2_B_writeaddr,
        dina      => IL_L1PHIE_PS10G_2_B_din,
        wea_out       => IL_L1PHIE_PS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIE_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIE_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIE_PS10G_2_B_start
      );

    IL_L1PHIF_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIF_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIF_PS10G_2_B_wea_delay,
        addra     => IL_L1PHIF_PS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIF_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIF_PS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIF_PS10G_2_B_V_dout,
        sync_nent => IL_L1PHIF_PS10G_2_B_start,
        nent_o    => IL_L1PHIF_PS10G_2_B_AV_dout_nent
      );

    IL_L1PHIF_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIF_PS10G_2_B_wea,
        addra     => IL_L1PHIF_PS10G_2_B_writeaddr,
        dina      => IL_L1PHIF_PS10G_2_B_din,
        wea_out       => IL_L1PHIF_PS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIF_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIF_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIF_PS10G_2_B_start
      );

    IL_L1PHIG_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIG_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIG_PS10G_2_B_wea_delay,
        addra     => IL_L1PHIG_PS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIG_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIG_PS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIG_PS10G_2_B_V_dout,
        sync_nent => IL_L1PHIG_PS10G_2_B_start,
        nent_o    => IL_L1PHIG_PS10G_2_B_AV_dout_nent
      );

    IL_L1PHIG_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIG_PS10G_2_B_wea,
        addra     => IL_L1PHIG_PS10G_2_B_writeaddr,
        dina      => IL_L1PHIG_PS10G_2_B_din,
        wea_out       => IL_L1PHIG_PS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIG_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIG_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIG_PS10G_2_B_start
      );

    IL_L1PHIH_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIH_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIH_PS10G_2_B_wea_delay,
        addra     => IL_L1PHIH_PS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIH_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIH_PS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIH_PS10G_2_B_V_dout,
        sync_nent => IL_L1PHIH_PS10G_2_B_start,
        nent_o    => IL_L1PHIH_PS10G_2_B_AV_dout_nent
      );

    IL_L1PHIH_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIH_PS10G_2_B_wea,
        addra     => IL_L1PHIH_PS10G_2_B_writeaddr,
        dina      => IL_L1PHIH_PS10G_2_B_din,
        wea_out       => IL_L1PHIH_PS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIH_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIH_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIH_PS10G_2_B_start
      );

    IL_D2PHIA_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_PS10G_2_A_wea_delay,
        addra     => IL_D2PHIA_PS10G_2_A_writeaddr_delay,
        dina      => IL_D2PHIA_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_PS10G_2_A_V_readaddr,
        doutb     => IL_D2PHIA_PS10G_2_A_V_dout,
        sync_nent => IL_D2PHIA_PS10G_2_A_start,
        nent_o    => IL_D2PHIA_PS10G_2_A_AV_dout_nent
      );

    IL_D2PHIA_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_PS10G_2_A_wea,
        addra     => IL_D2PHIA_PS10G_2_A_writeaddr,
        dina      => IL_D2PHIA_PS10G_2_A_din,
        wea_out       => IL_D2PHIA_PS10G_2_A_wea_delay,
        addra_out     => IL_D2PHIA_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_PS10G_2_A_start
      );

    IL_D2PHIB_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_PS10G_2_A_wea_delay,
        addra     => IL_D2PHIB_PS10G_2_A_writeaddr_delay,
        dina      => IL_D2PHIB_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_PS10G_2_A_V_readaddr,
        doutb     => IL_D2PHIB_PS10G_2_A_V_dout,
        sync_nent => IL_D2PHIB_PS10G_2_A_start,
        nent_o    => IL_D2PHIB_PS10G_2_A_AV_dout_nent
      );

    IL_D2PHIB_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_PS10G_2_A_wea,
        addra     => IL_D2PHIB_PS10G_2_A_writeaddr,
        dina      => IL_D2PHIB_PS10G_2_A_din,
        wea_out       => IL_D2PHIB_PS10G_2_A_wea_delay,
        addra_out     => IL_D2PHIB_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_PS10G_2_A_start
      );

    IL_D2PHIB_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_PS10G_2_B_wea_delay,
        addra     => IL_D2PHIB_PS10G_2_B_writeaddr_delay,
        dina      => IL_D2PHIB_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_PS10G_2_B_V_readaddr,
        doutb     => IL_D2PHIB_PS10G_2_B_V_dout,
        sync_nent => IL_D2PHIB_PS10G_2_B_start,
        nent_o    => IL_D2PHIB_PS10G_2_B_AV_dout_nent
      );

    IL_D2PHIB_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_PS10G_2_B_wea,
        addra     => IL_D2PHIB_PS10G_2_B_writeaddr,
        dina      => IL_D2PHIB_PS10G_2_B_din,
        wea_out       => IL_D2PHIB_PS10G_2_B_wea_delay,
        addra_out     => IL_D2PHIB_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_PS10G_2_B_start
      );

    IL_D2PHIC_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_PS10G_2_A_wea_delay,
        addra     => IL_D2PHIC_PS10G_2_A_writeaddr_delay,
        dina      => IL_D2PHIC_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_PS10G_2_A_V_readaddr,
        doutb     => IL_D2PHIC_PS10G_2_A_V_dout,
        sync_nent => IL_D2PHIC_PS10G_2_A_start,
        nent_o    => IL_D2PHIC_PS10G_2_A_AV_dout_nent
      );

    IL_D2PHIC_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_PS10G_2_A_wea,
        addra     => IL_D2PHIC_PS10G_2_A_writeaddr,
        dina      => IL_D2PHIC_PS10G_2_A_din,
        wea_out       => IL_D2PHIC_PS10G_2_A_wea_delay,
        addra_out     => IL_D2PHIC_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_PS10G_2_A_start
      );

    IL_D2PHIC_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_PS10G_2_B_wea_delay,
        addra     => IL_D2PHIC_PS10G_2_B_writeaddr_delay,
        dina      => IL_D2PHIC_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_PS10G_2_B_V_readaddr,
        doutb     => IL_D2PHIC_PS10G_2_B_V_dout,
        sync_nent => IL_D2PHIC_PS10G_2_B_start,
        nent_o    => IL_D2PHIC_PS10G_2_B_AV_dout_nent
      );

    IL_D2PHIC_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_PS10G_2_B_wea,
        addra     => IL_D2PHIC_PS10G_2_B_writeaddr,
        dina      => IL_D2PHIC_PS10G_2_B_din,
        wea_out       => IL_D2PHIC_PS10G_2_B_wea_delay,
        addra_out     => IL_D2PHIC_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_PS10G_2_B_start
      );

    IL_D2PHID_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_PS10G_2_B_wea_delay,
        addra     => IL_D2PHID_PS10G_2_B_writeaddr_delay,
        dina      => IL_D2PHID_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_PS10G_2_B_V_readaddr,
        doutb     => IL_D2PHID_PS10G_2_B_V_dout,
        sync_nent => IL_D2PHID_PS10G_2_B_start,
        nent_o    => IL_D2PHID_PS10G_2_B_AV_dout_nent
      );

    IL_D2PHID_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_PS10G_2_B_wea,
        addra     => IL_D2PHID_PS10G_2_B_writeaddr,
        dina      => IL_D2PHID_PS10G_2_B_din,
        wea_out       => IL_D2PHID_PS10G_2_B_wea_delay,
        addra_out     => IL_D2PHID_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_D2PHID_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_PS10G_2_B_start
      );

    IL_D4PHIA_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIA_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIA_PS10G_2_A_wea_delay,
        addra     => IL_D4PHIA_PS10G_2_A_writeaddr_delay,
        dina      => IL_D4PHIA_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIA_PS10G_2_A_V_readaddr,
        doutb     => IL_D4PHIA_PS10G_2_A_V_dout,
        sync_nent => IL_D4PHIA_PS10G_2_A_start,
        nent_o    => IL_D4PHIA_PS10G_2_A_AV_dout_nent
      );

    IL_D4PHIA_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIA_PS10G_2_A_wea,
        addra     => IL_D4PHIA_PS10G_2_A_writeaddr,
        dina      => IL_D4PHIA_PS10G_2_A_din,
        wea_out       => IL_D4PHIA_PS10G_2_A_wea_delay,
        addra_out     => IL_D4PHIA_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIA_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIA_PS10G_2_A_start
      );

    IL_D4PHIB_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_PS10G_2_A_wea_delay,
        addra     => IL_D4PHIB_PS10G_2_A_writeaddr_delay,
        dina      => IL_D4PHIB_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_PS10G_2_A_V_readaddr,
        doutb     => IL_D4PHIB_PS10G_2_A_V_dout,
        sync_nent => IL_D4PHIB_PS10G_2_A_start,
        nent_o    => IL_D4PHIB_PS10G_2_A_AV_dout_nent
      );

    IL_D4PHIB_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_PS10G_2_A_wea,
        addra     => IL_D4PHIB_PS10G_2_A_writeaddr,
        dina      => IL_D4PHIB_PS10G_2_A_din,
        wea_out       => IL_D4PHIB_PS10G_2_A_wea_delay,
        addra_out     => IL_D4PHIB_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIB_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_PS10G_2_A_start
      );

    IL_D4PHIB_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_PS10G_2_B_wea_delay,
        addra     => IL_D4PHIB_PS10G_2_B_writeaddr_delay,
        dina      => IL_D4PHIB_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_PS10G_2_B_V_readaddr,
        doutb     => IL_D4PHIB_PS10G_2_B_V_dout,
        sync_nent => IL_D4PHIB_PS10G_2_B_start,
        nent_o    => IL_D4PHIB_PS10G_2_B_AV_dout_nent
      );

    IL_D4PHIB_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_PS10G_2_B_wea,
        addra     => IL_D4PHIB_PS10G_2_B_writeaddr,
        dina      => IL_D4PHIB_PS10G_2_B_din,
        wea_out       => IL_D4PHIB_PS10G_2_B_wea_delay,
        addra_out     => IL_D4PHIB_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIB_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_PS10G_2_B_start
      );

    IL_D4PHIC_PS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_PS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_PS10G_2_A_wea_delay,
        addra     => IL_D4PHIC_PS10G_2_A_writeaddr_delay,
        dina      => IL_D4PHIC_PS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_PS10G_2_A_V_readaddr,
        doutb     => IL_D4PHIC_PS10G_2_A_V_dout,
        sync_nent => IL_D4PHIC_PS10G_2_A_start,
        nent_o    => IL_D4PHIC_PS10G_2_A_AV_dout_nent
      );

    IL_D4PHIC_PS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_PS10G_2_A_wea,
        addra     => IL_D4PHIC_PS10G_2_A_writeaddr,
        dina      => IL_D4PHIC_PS10G_2_A_din,
        wea_out       => IL_D4PHIC_PS10G_2_A_wea_delay,
        addra_out     => IL_D4PHIC_PS10G_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIC_PS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_PS10G_2_A_start
      );

    IL_D4PHIC_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_PS10G_2_B_wea_delay,
        addra     => IL_D4PHIC_PS10G_2_B_writeaddr_delay,
        dina      => IL_D4PHIC_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_PS10G_2_B_V_readaddr,
        doutb     => IL_D4PHIC_PS10G_2_B_V_dout,
        sync_nent => IL_D4PHIC_PS10G_2_B_start,
        nent_o    => IL_D4PHIC_PS10G_2_B_AV_dout_nent
      );

    IL_D4PHIC_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_PS10G_2_B_wea,
        addra     => IL_D4PHIC_PS10G_2_B_writeaddr,
        dina      => IL_D4PHIC_PS10G_2_B_din,
        wea_out       => IL_D4PHIC_PS10G_2_B_wea_delay,
        addra_out     => IL_D4PHIC_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIC_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_PS10G_2_B_start
      );

    IL_D4PHID_PS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHID_PS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHID_PS10G_2_B_wea_delay,
        addra     => IL_D4PHID_PS10G_2_B_writeaddr_delay,
        dina      => IL_D4PHID_PS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHID_PS10G_2_B_V_readaddr,
        doutb     => IL_D4PHID_PS10G_2_B_V_dout,
        sync_nent => IL_D4PHID_PS10G_2_B_start,
        nent_o    => IL_D4PHID_PS10G_2_B_AV_dout_nent
      );

    IL_D4PHID_PS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHID_PS10G_2_B_wea,
        addra     => IL_D4PHID_PS10G_2_B_writeaddr,
        dina      => IL_D4PHID_PS10G_2_B_din,
        wea_out       => IL_D4PHID_PS10G_2_B_wea_delay,
        addra_out     => IL_D4PHID_PS10G_2_B_writeaddr_delay,
        dina_out      => IL_D4PHID_PS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHID_PS10G_2_B_start
      );

    IL_L2PHIA_PS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIA_PS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIA_PS10G_3_A_wea_delay,
        addra     => IL_L2PHIA_PS10G_3_A_writeaddr_delay,
        dina      => IL_L2PHIA_PS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIA_PS10G_3_A_V_readaddr,
        doutb     => IL_L2PHIA_PS10G_3_A_V_dout,
        sync_nent => IL_L2PHIA_PS10G_3_A_start,
        nent_o    => IL_L2PHIA_PS10G_3_A_AV_dout_nent
      );

    IL_L2PHIA_PS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIA_PS10G_3_A_wea,
        addra     => IL_L2PHIA_PS10G_3_A_writeaddr,
        dina      => IL_L2PHIA_PS10G_3_A_din,
        wea_out       => IL_L2PHIA_PS10G_3_A_wea_delay,
        addra_out     => IL_L2PHIA_PS10G_3_A_writeaddr_delay,
        dina_out      => IL_L2PHIA_PS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_L2PHIA_PS10G_3_A_start
      );

    IL_L2PHIB_PS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIB_PS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIB_PS10G_3_A_wea_delay,
        addra     => IL_L2PHIB_PS10G_3_A_writeaddr_delay,
        dina      => IL_L2PHIB_PS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIB_PS10G_3_A_V_readaddr,
        doutb     => IL_L2PHIB_PS10G_3_A_V_dout,
        sync_nent => IL_L2PHIB_PS10G_3_A_start,
        nent_o    => IL_L2PHIB_PS10G_3_A_AV_dout_nent
      );

    IL_L2PHIB_PS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIB_PS10G_3_A_wea,
        addra     => IL_L2PHIB_PS10G_3_A_writeaddr,
        dina      => IL_L2PHIB_PS10G_3_A_din,
        wea_out       => IL_L2PHIB_PS10G_3_A_wea_delay,
        addra_out     => IL_L2PHIB_PS10G_3_A_writeaddr_delay,
        dina_out      => IL_L2PHIB_PS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_L2PHIB_PS10G_3_A_start
      );

    IL_L2PHIB_PS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIB_PS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIB_PS10G_3_B_wea_delay,
        addra     => IL_L2PHIB_PS10G_3_B_writeaddr_delay,
        dina      => IL_L2PHIB_PS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIB_PS10G_3_B_V_readaddr,
        doutb     => IL_L2PHIB_PS10G_3_B_V_dout,
        sync_nent => IL_L2PHIB_PS10G_3_B_start,
        nent_o    => IL_L2PHIB_PS10G_3_B_AV_dout_nent
      );

    IL_L2PHIB_PS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIB_PS10G_3_B_wea,
        addra     => IL_L2PHIB_PS10G_3_B_writeaddr,
        dina      => IL_L2PHIB_PS10G_3_B_din,
        wea_out       => IL_L2PHIB_PS10G_3_B_wea_delay,
        addra_out     => IL_L2PHIB_PS10G_3_B_writeaddr_delay,
        dina_out      => IL_L2PHIB_PS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_L2PHIB_PS10G_3_B_start
      );

    IL_L2PHIC_PS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIC_PS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIC_PS10G_3_A_wea_delay,
        addra     => IL_L2PHIC_PS10G_3_A_writeaddr_delay,
        dina      => IL_L2PHIC_PS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIC_PS10G_3_A_V_readaddr,
        doutb     => IL_L2PHIC_PS10G_3_A_V_dout,
        sync_nent => IL_L2PHIC_PS10G_3_A_start,
        nent_o    => IL_L2PHIC_PS10G_3_A_AV_dout_nent
      );

    IL_L2PHIC_PS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIC_PS10G_3_A_wea,
        addra     => IL_L2PHIC_PS10G_3_A_writeaddr,
        dina      => IL_L2PHIC_PS10G_3_A_din,
        wea_out       => IL_L2PHIC_PS10G_3_A_wea_delay,
        addra_out     => IL_L2PHIC_PS10G_3_A_writeaddr_delay,
        dina_out      => IL_L2PHIC_PS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_L2PHIC_PS10G_3_A_start
      );

    IL_L2PHIC_PS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIC_PS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIC_PS10G_3_B_wea_delay,
        addra     => IL_L2PHIC_PS10G_3_B_writeaddr_delay,
        dina      => IL_L2PHIC_PS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIC_PS10G_3_B_V_readaddr,
        doutb     => IL_L2PHIC_PS10G_3_B_V_dout,
        sync_nent => IL_L2PHIC_PS10G_3_B_start,
        nent_o    => IL_L2PHIC_PS10G_3_B_AV_dout_nent
      );

    IL_L2PHIC_PS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIC_PS10G_3_B_wea,
        addra     => IL_L2PHIC_PS10G_3_B_writeaddr,
        dina      => IL_L2PHIC_PS10G_3_B_din,
        wea_out       => IL_L2PHIC_PS10G_3_B_wea_delay,
        addra_out     => IL_L2PHIC_PS10G_3_B_writeaddr_delay,
        dina_out      => IL_L2PHIC_PS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_L2PHIC_PS10G_3_B_start
      );

    IL_L2PHID_PS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHID_PS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHID_PS10G_3_B_wea_delay,
        addra     => IL_L2PHID_PS10G_3_B_writeaddr_delay,
        dina      => IL_L2PHID_PS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHID_PS10G_3_B_V_readaddr,
        doutb     => IL_L2PHID_PS10G_3_B_V_dout,
        sync_nent => IL_L2PHID_PS10G_3_B_start,
        nent_o    => IL_L2PHID_PS10G_3_B_AV_dout_nent
      );

    IL_L2PHID_PS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHID_PS10G_3_B_wea,
        addra     => IL_L2PHID_PS10G_3_B_writeaddr,
        dina      => IL_L2PHID_PS10G_3_B_din,
        wea_out       => IL_L2PHID_PS10G_3_B_wea_delay,
        addra_out     => IL_L2PHID_PS10G_3_B_writeaddr_delay,
        dina_out      => IL_L2PHID_PS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_L2PHID_PS10G_3_B_start
      );

    IL_D2PHIA_PS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_PS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_PS10G_3_A_wea_delay,
        addra     => IL_D2PHIA_PS10G_3_A_writeaddr_delay,
        dina      => IL_D2PHIA_PS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_PS10G_3_A_V_readaddr,
        doutb     => IL_D2PHIA_PS10G_3_A_V_dout,
        sync_nent => IL_D2PHIA_PS10G_3_A_start,
        nent_o    => IL_D2PHIA_PS10G_3_A_AV_dout_nent
      );

    IL_D2PHIA_PS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_PS10G_3_A_wea,
        addra     => IL_D2PHIA_PS10G_3_A_writeaddr,
        dina      => IL_D2PHIA_PS10G_3_A_din,
        wea_out       => IL_D2PHIA_PS10G_3_A_wea_delay,
        addra_out     => IL_D2PHIA_PS10G_3_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_PS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_PS10G_3_A_start
      );

    IL_D2PHIB_PS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_PS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_PS10G_3_A_wea_delay,
        addra     => IL_D2PHIB_PS10G_3_A_writeaddr_delay,
        dina      => IL_D2PHIB_PS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_PS10G_3_A_V_readaddr,
        doutb     => IL_D2PHIB_PS10G_3_A_V_dout,
        sync_nent => IL_D2PHIB_PS10G_3_A_start,
        nent_o    => IL_D2PHIB_PS10G_3_A_AV_dout_nent
      );

    IL_D2PHIB_PS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_PS10G_3_A_wea,
        addra     => IL_D2PHIB_PS10G_3_A_writeaddr,
        dina      => IL_D2PHIB_PS10G_3_A_din,
        wea_out       => IL_D2PHIB_PS10G_3_A_wea_delay,
        addra_out     => IL_D2PHIB_PS10G_3_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_PS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_PS10G_3_A_start
      );

    IL_D2PHIB_PS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_PS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_PS10G_3_B_wea_delay,
        addra     => IL_D2PHIB_PS10G_3_B_writeaddr_delay,
        dina      => IL_D2PHIB_PS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_PS10G_3_B_V_readaddr,
        doutb     => IL_D2PHIB_PS10G_3_B_V_dout,
        sync_nent => IL_D2PHIB_PS10G_3_B_start,
        nent_o    => IL_D2PHIB_PS10G_3_B_AV_dout_nent
      );

    IL_D2PHIB_PS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_PS10G_3_B_wea,
        addra     => IL_D2PHIB_PS10G_3_B_writeaddr,
        dina      => IL_D2PHIB_PS10G_3_B_din,
        wea_out       => IL_D2PHIB_PS10G_3_B_wea_delay,
        addra_out     => IL_D2PHIB_PS10G_3_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_PS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_PS10G_3_B_start
      );

    IL_D2PHIC_PS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_PS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_PS10G_3_A_wea_delay,
        addra     => IL_D2PHIC_PS10G_3_A_writeaddr_delay,
        dina      => IL_D2PHIC_PS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_PS10G_3_A_V_readaddr,
        doutb     => IL_D2PHIC_PS10G_3_A_V_dout,
        sync_nent => IL_D2PHIC_PS10G_3_A_start,
        nent_o    => IL_D2PHIC_PS10G_3_A_AV_dout_nent
      );

    IL_D2PHIC_PS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_PS10G_3_A_wea,
        addra     => IL_D2PHIC_PS10G_3_A_writeaddr,
        dina      => IL_D2PHIC_PS10G_3_A_din,
        wea_out       => IL_D2PHIC_PS10G_3_A_wea_delay,
        addra_out     => IL_D2PHIC_PS10G_3_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_PS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_PS10G_3_A_start
      );

    IL_D2PHIC_PS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_PS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_PS10G_3_B_wea_delay,
        addra     => IL_D2PHIC_PS10G_3_B_writeaddr_delay,
        dina      => IL_D2PHIC_PS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_PS10G_3_B_V_readaddr,
        doutb     => IL_D2PHIC_PS10G_3_B_V_dout,
        sync_nent => IL_D2PHIC_PS10G_3_B_start,
        nent_o    => IL_D2PHIC_PS10G_3_B_AV_dout_nent
      );

    IL_D2PHIC_PS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_PS10G_3_B_wea,
        addra     => IL_D2PHIC_PS10G_3_B_writeaddr,
        dina      => IL_D2PHIC_PS10G_3_B_din,
        wea_out       => IL_D2PHIC_PS10G_3_B_wea_delay,
        addra_out     => IL_D2PHIC_PS10G_3_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_PS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_PS10G_3_B_start
      );

    IL_D2PHID_PS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_PS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_PS10G_3_B_wea_delay,
        addra     => IL_D2PHID_PS10G_3_B_writeaddr_delay,
        dina      => IL_D2PHID_PS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_PS10G_3_B_V_readaddr,
        doutb     => IL_D2PHID_PS10G_3_B_V_dout,
        sync_nent => IL_D2PHID_PS10G_3_B_start,
        nent_o    => IL_D2PHID_PS10G_3_B_AV_dout_nent
      );

    IL_D2PHID_PS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_PS10G_3_B_wea,
        addra     => IL_D2PHID_PS10G_3_B_writeaddr,
        dina      => IL_D2PHID_PS10G_3_B_din,
        wea_out       => IL_D2PHID_PS10G_3_B_wea_delay,
        addra_out     => IL_D2PHID_PS10G_3_B_writeaddr_delay,
        dina_out      => IL_D2PHID_PS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_PS10G_3_B_start
      );

    IL_D1PHIA_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIA_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIA_PS10G_4_A_wea_delay,
        addra     => IL_D1PHIA_PS10G_4_A_writeaddr_delay,
        dina      => IL_D1PHIA_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIA_PS10G_4_A_V_readaddr,
        doutb     => IL_D1PHIA_PS10G_4_A_V_dout,
        sync_nent => IL_D1PHIA_PS10G_4_A_start,
        nent_o    => IL_D1PHIA_PS10G_4_A_AV_dout_nent
      );

    IL_D1PHIA_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIA_PS10G_4_A_wea,
        addra     => IL_D1PHIA_PS10G_4_A_writeaddr,
        dina      => IL_D1PHIA_PS10G_4_A_din,
        wea_out       => IL_D1PHIA_PS10G_4_A_wea_delay,
        addra_out     => IL_D1PHIA_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D1PHIA_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIA_PS10G_4_A_start
      );

    IL_D1PHIB_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_PS10G_4_A_wea_delay,
        addra     => IL_D1PHIB_PS10G_4_A_writeaddr_delay,
        dina      => IL_D1PHIB_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_PS10G_4_A_V_readaddr,
        doutb     => IL_D1PHIB_PS10G_4_A_V_dout,
        sync_nent => IL_D1PHIB_PS10G_4_A_start,
        nent_o    => IL_D1PHIB_PS10G_4_A_AV_dout_nent
      );

    IL_D1PHIB_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_PS10G_4_A_wea,
        addra     => IL_D1PHIB_PS10G_4_A_writeaddr,
        dina      => IL_D1PHIB_PS10G_4_A_din,
        wea_out       => IL_D1PHIB_PS10G_4_A_wea_delay,
        addra_out     => IL_D1PHIB_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D1PHIB_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_PS10G_4_A_start
      );

    IL_D1PHIB_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_PS10G_4_B_wea_delay,
        addra     => IL_D1PHIB_PS10G_4_B_writeaddr_delay,
        dina      => IL_D1PHIB_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_PS10G_4_B_V_readaddr,
        doutb     => IL_D1PHIB_PS10G_4_B_V_dout,
        sync_nent => IL_D1PHIB_PS10G_4_B_start,
        nent_o    => IL_D1PHIB_PS10G_4_B_AV_dout_nent
      );

    IL_D1PHIB_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_PS10G_4_B_wea,
        addra     => IL_D1PHIB_PS10G_4_B_writeaddr,
        dina      => IL_D1PHIB_PS10G_4_B_din,
        wea_out       => IL_D1PHIB_PS10G_4_B_wea_delay,
        addra_out     => IL_D1PHIB_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D1PHIB_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_PS10G_4_B_start
      );

    IL_D1PHIC_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_PS10G_4_A_wea_delay,
        addra     => IL_D1PHIC_PS10G_4_A_writeaddr_delay,
        dina      => IL_D1PHIC_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_PS10G_4_A_V_readaddr,
        doutb     => IL_D1PHIC_PS10G_4_A_V_dout,
        sync_nent => IL_D1PHIC_PS10G_4_A_start,
        nent_o    => IL_D1PHIC_PS10G_4_A_AV_dout_nent
      );

    IL_D1PHIC_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_PS10G_4_A_wea,
        addra     => IL_D1PHIC_PS10G_4_A_writeaddr,
        dina      => IL_D1PHIC_PS10G_4_A_din,
        wea_out       => IL_D1PHIC_PS10G_4_A_wea_delay,
        addra_out     => IL_D1PHIC_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D1PHIC_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_PS10G_4_A_start
      );

    IL_D1PHIC_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_PS10G_4_B_wea_delay,
        addra     => IL_D1PHIC_PS10G_4_B_writeaddr_delay,
        dina      => IL_D1PHIC_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_PS10G_4_B_V_readaddr,
        doutb     => IL_D1PHIC_PS10G_4_B_V_dout,
        sync_nent => IL_D1PHIC_PS10G_4_B_start,
        nent_o    => IL_D1PHIC_PS10G_4_B_AV_dout_nent
      );

    IL_D1PHIC_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_PS10G_4_B_wea,
        addra     => IL_D1PHIC_PS10G_4_B_writeaddr,
        dina      => IL_D1PHIC_PS10G_4_B_din,
        wea_out       => IL_D1PHIC_PS10G_4_B_wea_delay,
        addra_out     => IL_D1PHIC_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D1PHIC_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_PS10G_4_B_start
      );

    IL_D1PHID_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHID_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHID_PS10G_4_B_wea_delay,
        addra     => IL_D1PHID_PS10G_4_B_writeaddr_delay,
        dina      => IL_D1PHID_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHID_PS10G_4_B_V_readaddr,
        doutb     => IL_D1PHID_PS10G_4_B_V_dout,
        sync_nent => IL_D1PHID_PS10G_4_B_start,
        nent_o    => IL_D1PHID_PS10G_4_B_AV_dout_nent
      );

    IL_D1PHID_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHID_PS10G_4_B_wea,
        addra     => IL_D1PHID_PS10G_4_B_writeaddr,
        dina      => IL_D1PHID_PS10G_4_B_din,
        wea_out       => IL_D1PHID_PS10G_4_B_wea_delay,
        addra_out     => IL_D1PHID_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D1PHID_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHID_PS10G_4_B_start
      );

    IL_D3PHIA_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIA_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIA_PS10G_4_A_wea_delay,
        addra     => IL_D3PHIA_PS10G_4_A_writeaddr_delay,
        dina      => IL_D3PHIA_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIA_PS10G_4_A_V_readaddr,
        doutb     => IL_D3PHIA_PS10G_4_A_V_dout,
        sync_nent => IL_D3PHIA_PS10G_4_A_start,
        nent_o    => IL_D3PHIA_PS10G_4_A_AV_dout_nent
      );

    IL_D3PHIA_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIA_PS10G_4_A_wea,
        addra     => IL_D3PHIA_PS10G_4_A_writeaddr,
        dina      => IL_D3PHIA_PS10G_4_A_din,
        wea_out       => IL_D3PHIA_PS10G_4_A_wea_delay,
        addra_out     => IL_D3PHIA_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIA_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIA_PS10G_4_A_start
      );

    IL_D3PHIB_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_PS10G_4_A_wea_delay,
        addra     => IL_D3PHIB_PS10G_4_A_writeaddr_delay,
        dina      => IL_D3PHIB_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_PS10G_4_A_V_readaddr,
        doutb     => IL_D3PHIB_PS10G_4_A_V_dout,
        sync_nent => IL_D3PHIB_PS10G_4_A_start,
        nent_o    => IL_D3PHIB_PS10G_4_A_AV_dout_nent
      );

    IL_D3PHIB_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_PS10G_4_A_wea,
        addra     => IL_D3PHIB_PS10G_4_A_writeaddr,
        dina      => IL_D3PHIB_PS10G_4_A_din,
        wea_out       => IL_D3PHIB_PS10G_4_A_wea_delay,
        addra_out     => IL_D3PHIB_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIB_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_PS10G_4_A_start
      );

    IL_D3PHIB_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_PS10G_4_B_wea_delay,
        addra     => IL_D3PHIB_PS10G_4_B_writeaddr_delay,
        dina      => IL_D3PHIB_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_PS10G_4_B_V_readaddr,
        doutb     => IL_D3PHIB_PS10G_4_B_V_dout,
        sync_nent => IL_D3PHIB_PS10G_4_B_start,
        nent_o    => IL_D3PHIB_PS10G_4_B_AV_dout_nent
      );

    IL_D3PHIB_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_PS10G_4_B_wea,
        addra     => IL_D3PHIB_PS10G_4_B_writeaddr,
        dina      => IL_D3PHIB_PS10G_4_B_din,
        wea_out       => IL_D3PHIB_PS10G_4_B_wea_delay,
        addra_out     => IL_D3PHIB_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIB_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_PS10G_4_B_start
      );

    IL_D3PHIC_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_PS10G_4_A_wea_delay,
        addra     => IL_D3PHIC_PS10G_4_A_writeaddr_delay,
        dina      => IL_D3PHIC_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_PS10G_4_A_V_readaddr,
        doutb     => IL_D3PHIC_PS10G_4_A_V_dout,
        sync_nent => IL_D3PHIC_PS10G_4_A_start,
        nent_o    => IL_D3PHIC_PS10G_4_A_AV_dout_nent
      );

    IL_D3PHIC_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_PS10G_4_A_wea,
        addra     => IL_D3PHIC_PS10G_4_A_writeaddr,
        dina      => IL_D3PHIC_PS10G_4_A_din,
        wea_out       => IL_D3PHIC_PS10G_4_A_wea_delay,
        addra_out     => IL_D3PHIC_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIC_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_PS10G_4_A_start
      );

    IL_D3PHIC_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_PS10G_4_B_wea_delay,
        addra     => IL_D3PHIC_PS10G_4_B_writeaddr_delay,
        dina      => IL_D3PHIC_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_PS10G_4_B_V_readaddr,
        doutb     => IL_D3PHIC_PS10G_4_B_V_dout,
        sync_nent => IL_D3PHIC_PS10G_4_B_start,
        nent_o    => IL_D3PHIC_PS10G_4_B_AV_dout_nent
      );

    IL_D3PHIC_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_PS10G_4_B_wea,
        addra     => IL_D3PHIC_PS10G_4_B_writeaddr,
        dina      => IL_D3PHIC_PS10G_4_B_din,
        wea_out       => IL_D3PHIC_PS10G_4_B_wea_delay,
        addra_out     => IL_D3PHIC_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIC_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_PS10G_4_B_start
      );

    IL_D3PHID_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHID_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHID_PS10G_4_B_wea_delay,
        addra     => IL_D3PHID_PS10G_4_B_writeaddr_delay,
        dina      => IL_D3PHID_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHID_PS10G_4_B_V_readaddr,
        doutb     => IL_D3PHID_PS10G_4_B_V_dout,
        sync_nent => IL_D3PHID_PS10G_4_B_start,
        nent_o    => IL_D3PHID_PS10G_4_B_AV_dout_nent
      );

    IL_D3PHID_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHID_PS10G_4_B_wea,
        addra     => IL_D3PHID_PS10G_4_B_writeaddr,
        dina      => IL_D3PHID_PS10G_4_B_din,
        wea_out       => IL_D3PHID_PS10G_4_B_wea_delay,
        addra_out     => IL_D3PHID_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D3PHID_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHID_PS10G_4_B_start
      );

    IL_D5PHIA_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIA_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIA_PS10G_4_A_wea_delay,
        addra     => IL_D5PHIA_PS10G_4_A_writeaddr_delay,
        dina      => IL_D5PHIA_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIA_PS10G_4_A_V_readaddr,
        doutb     => IL_D5PHIA_PS10G_4_A_V_dout,
        sync_nent => IL_D5PHIA_PS10G_4_A_start,
        nent_o    => IL_D5PHIA_PS10G_4_A_AV_dout_nent
      );

    IL_D5PHIA_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIA_PS10G_4_A_wea,
        addra     => IL_D5PHIA_PS10G_4_A_writeaddr,
        dina      => IL_D5PHIA_PS10G_4_A_din,
        wea_out       => IL_D5PHIA_PS10G_4_A_wea_delay,
        addra_out     => IL_D5PHIA_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D5PHIA_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIA_PS10G_4_A_start
      );

    IL_D5PHIB_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_PS10G_4_A_wea_delay,
        addra     => IL_D5PHIB_PS10G_4_A_writeaddr_delay,
        dina      => IL_D5PHIB_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_PS10G_4_A_V_readaddr,
        doutb     => IL_D5PHIB_PS10G_4_A_V_dout,
        sync_nent => IL_D5PHIB_PS10G_4_A_start,
        nent_o    => IL_D5PHIB_PS10G_4_A_AV_dout_nent
      );

    IL_D5PHIB_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_PS10G_4_A_wea,
        addra     => IL_D5PHIB_PS10G_4_A_writeaddr,
        dina      => IL_D5PHIB_PS10G_4_A_din,
        wea_out       => IL_D5PHIB_PS10G_4_A_wea_delay,
        addra_out     => IL_D5PHIB_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D5PHIB_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_PS10G_4_A_start
      );

    IL_D5PHIB_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_PS10G_4_B_wea_delay,
        addra     => IL_D5PHIB_PS10G_4_B_writeaddr_delay,
        dina      => IL_D5PHIB_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_PS10G_4_B_V_readaddr,
        doutb     => IL_D5PHIB_PS10G_4_B_V_dout,
        sync_nent => IL_D5PHIB_PS10G_4_B_start,
        nent_o    => IL_D5PHIB_PS10G_4_B_AV_dout_nent
      );

    IL_D5PHIB_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_PS10G_4_B_wea,
        addra     => IL_D5PHIB_PS10G_4_B_writeaddr,
        dina      => IL_D5PHIB_PS10G_4_B_din,
        wea_out       => IL_D5PHIB_PS10G_4_B_wea_delay,
        addra_out     => IL_D5PHIB_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D5PHIB_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_PS10G_4_B_start
      );

    IL_D5PHIC_PS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_PS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_PS10G_4_A_wea_delay,
        addra     => IL_D5PHIC_PS10G_4_A_writeaddr_delay,
        dina      => IL_D5PHIC_PS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_PS10G_4_A_V_readaddr,
        doutb     => IL_D5PHIC_PS10G_4_A_V_dout,
        sync_nent => IL_D5PHIC_PS10G_4_A_start,
        nent_o    => IL_D5PHIC_PS10G_4_A_AV_dout_nent
      );

    IL_D5PHIC_PS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_PS10G_4_A_wea,
        addra     => IL_D5PHIC_PS10G_4_A_writeaddr,
        dina      => IL_D5PHIC_PS10G_4_A_din,
        wea_out       => IL_D5PHIC_PS10G_4_A_wea_delay,
        addra_out     => IL_D5PHIC_PS10G_4_A_writeaddr_delay,
        dina_out      => IL_D5PHIC_PS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_PS10G_4_A_start
      );

    IL_D5PHIC_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_PS10G_4_B_wea_delay,
        addra     => IL_D5PHIC_PS10G_4_B_writeaddr_delay,
        dina      => IL_D5PHIC_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_PS10G_4_B_V_readaddr,
        doutb     => IL_D5PHIC_PS10G_4_B_V_dout,
        sync_nent => IL_D5PHIC_PS10G_4_B_start,
        nent_o    => IL_D5PHIC_PS10G_4_B_AV_dout_nent
      );

    IL_D5PHIC_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_PS10G_4_B_wea,
        addra     => IL_D5PHIC_PS10G_4_B_writeaddr,
        dina      => IL_D5PHIC_PS10G_4_B_din,
        wea_out       => IL_D5PHIC_PS10G_4_B_wea_delay,
        addra_out     => IL_D5PHIC_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D5PHIC_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_PS10G_4_B_start
      );

    IL_D5PHID_PS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHID_PS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHID_PS10G_4_B_wea_delay,
        addra     => IL_D5PHID_PS10G_4_B_writeaddr_delay,
        dina      => IL_D5PHID_PS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHID_PS10G_4_B_V_readaddr,
        doutb     => IL_D5PHID_PS10G_4_B_V_dout,
        sync_nent => IL_D5PHID_PS10G_4_B_start,
        nent_o    => IL_D5PHID_PS10G_4_B_AV_dout_nent
      );

    IL_D5PHID_PS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHID_PS10G_4_B_wea,
        addra     => IL_D5PHID_PS10G_4_B_writeaddr,
        dina      => IL_D5PHID_PS10G_4_B_din,
        wea_out       => IL_D5PHID_PS10G_4_B_wea_delay,
        addra_out     => IL_D5PHID_PS10G_4_B_writeaddr_delay,
        dina_out      => IL_D5PHID_PS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHID_PS10G_4_B_start
      );

    IL_L3PHIA_PS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIA_PS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIA_PS_1_A_wea_delay,
        addra     => IL_L3PHIA_PS_1_A_writeaddr_delay,
        dina      => IL_L3PHIA_PS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIA_PS_1_A_V_readaddr,
        doutb     => IL_L3PHIA_PS_1_A_V_dout,
        sync_nent => IL_L3PHIA_PS_1_A_start,
        nent_o    => IL_L3PHIA_PS_1_A_AV_dout_nent
      );

    IL_L3PHIA_PS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIA_PS_1_A_wea,
        addra     => IL_L3PHIA_PS_1_A_writeaddr,
        dina      => IL_L3PHIA_PS_1_A_din,
        wea_out       => IL_L3PHIA_PS_1_A_wea_delay,
        addra_out     => IL_L3PHIA_PS_1_A_writeaddr_delay,
        dina_out      => IL_L3PHIA_PS_1_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIA_PS_1_A_start
      );

    IL_L3PHIB_PS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIB_PS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIB_PS_1_A_wea_delay,
        addra     => IL_L3PHIB_PS_1_A_writeaddr_delay,
        dina      => IL_L3PHIB_PS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIB_PS_1_A_V_readaddr,
        doutb     => IL_L3PHIB_PS_1_A_V_dout,
        sync_nent => IL_L3PHIB_PS_1_A_start,
        nent_o    => IL_L3PHIB_PS_1_A_AV_dout_nent
      );

    IL_L3PHIB_PS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIB_PS_1_A_wea,
        addra     => IL_L3PHIB_PS_1_A_writeaddr,
        dina      => IL_L3PHIB_PS_1_A_din,
        wea_out       => IL_L3PHIB_PS_1_A_wea_delay,
        addra_out     => IL_L3PHIB_PS_1_A_writeaddr_delay,
        dina_out      => IL_L3PHIB_PS_1_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIB_PS_1_A_start
      );

    IL_L3PHIC_PS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIC_PS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIC_PS_1_B_wea_delay,
        addra     => IL_L3PHIC_PS_1_B_writeaddr_delay,
        dina      => IL_L3PHIC_PS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIC_PS_1_B_V_readaddr,
        doutb     => IL_L3PHIC_PS_1_B_V_dout,
        sync_nent => IL_L3PHIC_PS_1_B_start,
        nent_o    => IL_L3PHIC_PS_1_B_AV_dout_nent
      );

    IL_L3PHIC_PS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIC_PS_1_B_wea,
        addra     => IL_L3PHIC_PS_1_B_writeaddr,
        dina      => IL_L3PHIC_PS_1_B_din,
        wea_out       => IL_L3PHIC_PS_1_B_wea_delay,
        addra_out     => IL_L3PHIC_PS_1_B_writeaddr_delay,
        dina_out      => IL_L3PHIC_PS_1_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHIC_PS_1_B_start
      );

    IL_L3PHID_PS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHID_PS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHID_PS_1_B_wea_delay,
        addra     => IL_L3PHID_PS_1_B_writeaddr_delay,
        dina      => IL_L3PHID_PS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHID_PS_1_B_V_readaddr,
        doutb     => IL_L3PHID_PS_1_B_V_dout,
        sync_nent => IL_L3PHID_PS_1_B_start,
        nent_o    => IL_L3PHID_PS_1_B_AV_dout_nent
      );

    IL_L3PHID_PS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHID_PS_1_B_wea,
        addra     => IL_L3PHID_PS_1_B_writeaddr,
        dina      => IL_L3PHID_PS_1_B_din,
        wea_out       => IL_L3PHID_PS_1_B_wea_delay,
        addra_out     => IL_L3PHID_PS_1_B_writeaddr_delay,
        dina_out      => IL_L3PHID_PS_1_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHID_PS_1_B_start
      );

    IL_D2PHIA_PS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_PS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_PS_1_A_wea_delay,
        addra     => IL_D2PHIA_PS_1_A_writeaddr_delay,
        dina      => IL_D2PHIA_PS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_PS_1_A_V_readaddr,
        doutb     => IL_D2PHIA_PS_1_A_V_dout,
        sync_nent => IL_D2PHIA_PS_1_A_start,
        nent_o    => IL_D2PHIA_PS_1_A_AV_dout_nent
      );

    IL_D2PHIA_PS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_PS_1_A_wea,
        addra     => IL_D2PHIA_PS_1_A_writeaddr,
        dina      => IL_D2PHIA_PS_1_A_din,
        wea_out       => IL_D2PHIA_PS_1_A_wea_delay,
        addra_out     => IL_D2PHIA_PS_1_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_PS_1_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_PS_1_A_start
      );

    IL_D2PHIB_PS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_PS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_PS_1_A_wea_delay,
        addra     => IL_D2PHIB_PS_1_A_writeaddr_delay,
        dina      => IL_D2PHIB_PS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_PS_1_A_V_readaddr,
        doutb     => IL_D2PHIB_PS_1_A_V_dout,
        sync_nent => IL_D2PHIB_PS_1_A_start,
        nent_o    => IL_D2PHIB_PS_1_A_AV_dout_nent
      );

    IL_D2PHIB_PS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_PS_1_A_wea,
        addra     => IL_D2PHIB_PS_1_A_writeaddr,
        dina      => IL_D2PHIB_PS_1_A_din,
        wea_out       => IL_D2PHIB_PS_1_A_wea_delay,
        addra_out     => IL_D2PHIB_PS_1_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_PS_1_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_PS_1_A_start
      );

    IL_D2PHIB_PS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_PS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_PS_1_B_wea_delay,
        addra     => IL_D2PHIB_PS_1_B_writeaddr_delay,
        dina      => IL_D2PHIB_PS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_PS_1_B_V_readaddr,
        doutb     => IL_D2PHIB_PS_1_B_V_dout,
        sync_nent => IL_D2PHIB_PS_1_B_start,
        nent_o    => IL_D2PHIB_PS_1_B_AV_dout_nent
      );

    IL_D2PHIB_PS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_PS_1_B_wea,
        addra     => IL_D2PHIB_PS_1_B_writeaddr,
        dina      => IL_D2PHIB_PS_1_B_din,
        wea_out       => IL_D2PHIB_PS_1_B_wea_delay,
        addra_out     => IL_D2PHIB_PS_1_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_PS_1_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_PS_1_B_start
      );

    IL_D2PHIC_PS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_PS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_PS_1_A_wea_delay,
        addra     => IL_D2PHIC_PS_1_A_writeaddr_delay,
        dina      => IL_D2PHIC_PS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_PS_1_A_V_readaddr,
        doutb     => IL_D2PHIC_PS_1_A_V_dout,
        sync_nent => IL_D2PHIC_PS_1_A_start,
        nent_o    => IL_D2PHIC_PS_1_A_AV_dout_nent
      );

    IL_D2PHIC_PS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_PS_1_A_wea,
        addra     => IL_D2PHIC_PS_1_A_writeaddr,
        dina      => IL_D2PHIC_PS_1_A_din,
        wea_out       => IL_D2PHIC_PS_1_A_wea_delay,
        addra_out     => IL_D2PHIC_PS_1_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_PS_1_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_PS_1_A_start
      );

    IL_D2PHIC_PS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_PS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_PS_1_B_wea_delay,
        addra     => IL_D2PHIC_PS_1_B_writeaddr_delay,
        dina      => IL_D2PHIC_PS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_PS_1_B_V_readaddr,
        doutb     => IL_D2PHIC_PS_1_B_V_dout,
        sync_nent => IL_D2PHIC_PS_1_B_start,
        nent_o    => IL_D2PHIC_PS_1_B_AV_dout_nent
      );

    IL_D2PHIC_PS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_PS_1_B_wea,
        addra     => IL_D2PHIC_PS_1_B_writeaddr,
        dina      => IL_D2PHIC_PS_1_B_din,
        wea_out       => IL_D2PHIC_PS_1_B_wea_delay,
        addra_out     => IL_D2PHIC_PS_1_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_PS_1_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_PS_1_B_start
      );

    IL_D2PHID_PS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_PS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_PS_1_B_wea_delay,
        addra     => IL_D2PHID_PS_1_B_writeaddr_delay,
        dina      => IL_D2PHID_PS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_PS_1_B_V_readaddr,
        doutb     => IL_D2PHID_PS_1_B_V_dout,
        sync_nent => IL_D2PHID_PS_1_B_start,
        nent_o    => IL_D2PHID_PS_1_B_AV_dout_nent
      );

    IL_D2PHID_PS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_PS_1_B_wea,
        addra     => IL_D2PHID_PS_1_B_writeaddr,
        dina      => IL_D2PHID_PS_1_B_din,
        wea_out       => IL_D2PHID_PS_1_B_wea_delay,
        addra_out     => IL_D2PHID_PS_1_B_writeaddr_delay,
        dina_out      => IL_D2PHID_PS_1_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_PS_1_B_start
      );

    IL_L3PHIA_PS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIA_PS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIA_PS_2_A_wea_delay,
        addra     => IL_L3PHIA_PS_2_A_writeaddr_delay,
        dina      => IL_L3PHIA_PS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIA_PS_2_A_V_readaddr,
        doutb     => IL_L3PHIA_PS_2_A_V_dout,
        sync_nent => IL_L3PHIA_PS_2_A_start,
        nent_o    => IL_L3PHIA_PS_2_A_AV_dout_nent
      );

    IL_L3PHIA_PS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIA_PS_2_A_wea,
        addra     => IL_L3PHIA_PS_2_A_writeaddr,
        dina      => IL_L3PHIA_PS_2_A_din,
        wea_out       => IL_L3PHIA_PS_2_A_wea_delay,
        addra_out     => IL_L3PHIA_PS_2_A_writeaddr_delay,
        dina_out      => IL_L3PHIA_PS_2_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIA_PS_2_A_start
      );

    IL_L3PHIB_PS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIB_PS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIB_PS_2_A_wea_delay,
        addra     => IL_L3PHIB_PS_2_A_writeaddr_delay,
        dina      => IL_L3PHIB_PS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIB_PS_2_A_V_readaddr,
        doutb     => IL_L3PHIB_PS_2_A_V_dout,
        sync_nent => IL_L3PHIB_PS_2_A_start,
        nent_o    => IL_L3PHIB_PS_2_A_AV_dout_nent
      );

    IL_L3PHIB_PS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIB_PS_2_A_wea,
        addra     => IL_L3PHIB_PS_2_A_writeaddr,
        dina      => IL_L3PHIB_PS_2_A_din,
        wea_out       => IL_L3PHIB_PS_2_A_wea_delay,
        addra_out     => IL_L3PHIB_PS_2_A_writeaddr_delay,
        dina_out      => IL_L3PHIB_PS_2_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIB_PS_2_A_start
      );

    IL_L3PHIB_PS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIB_PS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIB_PS_2_B_wea_delay,
        addra     => IL_L3PHIB_PS_2_B_writeaddr_delay,
        dina      => IL_L3PHIB_PS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIB_PS_2_B_V_readaddr,
        doutb     => IL_L3PHIB_PS_2_B_V_dout,
        sync_nent => IL_L3PHIB_PS_2_B_start,
        nent_o    => IL_L3PHIB_PS_2_B_AV_dout_nent
      );

    IL_L3PHIB_PS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIB_PS_2_B_wea,
        addra     => IL_L3PHIB_PS_2_B_writeaddr,
        dina      => IL_L3PHIB_PS_2_B_din,
        wea_out       => IL_L3PHIB_PS_2_B_wea_delay,
        addra_out     => IL_L3PHIB_PS_2_B_writeaddr_delay,
        dina_out      => IL_L3PHIB_PS_2_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHIB_PS_2_B_start
      );

    IL_L3PHIC_PS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIC_PS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIC_PS_2_B_wea_delay,
        addra     => IL_L3PHIC_PS_2_B_writeaddr_delay,
        dina      => IL_L3PHIC_PS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIC_PS_2_B_V_readaddr,
        doutb     => IL_L3PHIC_PS_2_B_V_dout,
        sync_nent => IL_L3PHIC_PS_2_B_start,
        nent_o    => IL_L3PHIC_PS_2_B_AV_dout_nent
      );

    IL_L3PHIC_PS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIC_PS_2_B_wea,
        addra     => IL_L3PHIC_PS_2_B_writeaddr,
        dina      => IL_L3PHIC_PS_2_B_din,
        wea_out       => IL_L3PHIC_PS_2_B_wea_delay,
        addra_out     => IL_L3PHIC_PS_2_B_writeaddr_delay,
        dina_out      => IL_L3PHIC_PS_2_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHIC_PS_2_B_start
      );

    IL_L3PHID_PS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHID_PS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHID_PS_2_B_wea_delay,
        addra     => IL_L3PHID_PS_2_B_writeaddr_delay,
        dina      => IL_L3PHID_PS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHID_PS_2_B_V_readaddr,
        doutb     => IL_L3PHID_PS_2_B_V_dout,
        sync_nent => IL_L3PHID_PS_2_B_start,
        nent_o    => IL_L3PHID_PS_2_B_AV_dout_nent
      );

    IL_L3PHID_PS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHID_PS_2_B_wea,
        addra     => IL_L3PHID_PS_2_B_writeaddr,
        dina      => IL_L3PHID_PS_2_B_din,
        wea_out       => IL_L3PHID_PS_2_B_wea_delay,
        addra_out     => IL_L3PHID_PS_2_B_writeaddr_delay,
        dina_out      => IL_L3PHID_PS_2_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHID_PS_2_B_start
      );

    IL_D4PHIA_PS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIA_PS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIA_PS_2_A_wea_delay,
        addra     => IL_D4PHIA_PS_2_A_writeaddr_delay,
        dina      => IL_D4PHIA_PS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIA_PS_2_A_V_readaddr,
        doutb     => IL_D4PHIA_PS_2_A_V_dout,
        sync_nent => IL_D4PHIA_PS_2_A_start,
        nent_o    => IL_D4PHIA_PS_2_A_AV_dout_nent
      );

    IL_D4PHIA_PS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIA_PS_2_A_wea,
        addra     => IL_D4PHIA_PS_2_A_writeaddr,
        dina      => IL_D4PHIA_PS_2_A_din,
        wea_out       => IL_D4PHIA_PS_2_A_wea_delay,
        addra_out     => IL_D4PHIA_PS_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIA_PS_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIA_PS_2_A_start
      );

    IL_D4PHIB_PS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_PS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_PS_2_A_wea_delay,
        addra     => IL_D4PHIB_PS_2_A_writeaddr_delay,
        dina      => IL_D4PHIB_PS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_PS_2_A_V_readaddr,
        doutb     => IL_D4PHIB_PS_2_A_V_dout,
        sync_nent => IL_D4PHIB_PS_2_A_start,
        nent_o    => IL_D4PHIB_PS_2_A_AV_dout_nent
      );

    IL_D4PHIB_PS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_PS_2_A_wea,
        addra     => IL_D4PHIB_PS_2_A_writeaddr,
        dina      => IL_D4PHIB_PS_2_A_din,
        wea_out       => IL_D4PHIB_PS_2_A_wea_delay,
        addra_out     => IL_D4PHIB_PS_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIB_PS_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_PS_2_A_start
      );

    IL_D4PHIB_PS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_PS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_PS_2_B_wea_delay,
        addra     => IL_D4PHIB_PS_2_B_writeaddr_delay,
        dina      => IL_D4PHIB_PS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_PS_2_B_V_readaddr,
        doutb     => IL_D4PHIB_PS_2_B_V_dout,
        sync_nent => IL_D4PHIB_PS_2_B_start,
        nent_o    => IL_D4PHIB_PS_2_B_AV_dout_nent
      );

    IL_D4PHIB_PS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_PS_2_B_wea,
        addra     => IL_D4PHIB_PS_2_B_writeaddr,
        dina      => IL_D4PHIB_PS_2_B_din,
        wea_out       => IL_D4PHIB_PS_2_B_wea_delay,
        addra_out     => IL_D4PHIB_PS_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIB_PS_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_PS_2_B_start
      );

    IL_D4PHIC_PS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_PS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_PS_2_A_wea_delay,
        addra     => IL_D4PHIC_PS_2_A_writeaddr_delay,
        dina      => IL_D4PHIC_PS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_PS_2_A_V_readaddr,
        doutb     => IL_D4PHIC_PS_2_A_V_dout,
        sync_nent => IL_D4PHIC_PS_2_A_start,
        nent_o    => IL_D4PHIC_PS_2_A_AV_dout_nent
      );

    IL_D4PHIC_PS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_PS_2_A_wea,
        addra     => IL_D4PHIC_PS_2_A_writeaddr,
        dina      => IL_D4PHIC_PS_2_A_din,
        wea_out       => IL_D4PHIC_PS_2_A_wea_delay,
        addra_out     => IL_D4PHIC_PS_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIC_PS_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_PS_2_A_start
      );

    IL_D4PHIC_PS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_PS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_PS_2_B_wea_delay,
        addra     => IL_D4PHIC_PS_2_B_writeaddr_delay,
        dina      => IL_D4PHIC_PS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_PS_2_B_V_readaddr,
        doutb     => IL_D4PHIC_PS_2_B_V_dout,
        sync_nent => IL_D4PHIC_PS_2_B_start,
        nent_o    => IL_D4PHIC_PS_2_B_AV_dout_nent
      );

    IL_D4PHIC_PS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_PS_2_B_wea,
        addra     => IL_D4PHIC_PS_2_B_writeaddr,
        dina      => IL_D4PHIC_PS_2_B_din,
        wea_out       => IL_D4PHIC_PS_2_B_wea_delay,
        addra_out     => IL_D4PHIC_PS_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIC_PS_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_PS_2_B_start
      );

    IL_D4PHID_PS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHID_PS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHID_PS_2_B_wea_delay,
        addra     => IL_D4PHID_PS_2_B_writeaddr_delay,
        dina      => IL_D4PHID_PS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHID_PS_2_B_V_readaddr,
        doutb     => IL_D4PHID_PS_2_B_V_dout,
        sync_nent => IL_D4PHID_PS_2_B_start,
        nent_o    => IL_D4PHID_PS_2_B_AV_dout_nent
      );

    IL_D4PHID_PS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHID_PS_2_B_wea,
        addra     => IL_D4PHID_PS_2_B_writeaddr,
        dina      => IL_D4PHID_PS_2_B_din,
        wea_out       => IL_D4PHID_PS_2_B_wea_delay,
        addra_out     => IL_D4PHID_PS_2_B_writeaddr_delay,
        dina_out      => IL_D4PHID_PS_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHID_PS_2_B_start
      );

    IL_L1PHIA_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIA_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIA_negPS10G_1_A_wea_delay,
        addra     => IL_L1PHIA_negPS10G_1_A_writeaddr_delay,
        dina      => IL_L1PHIA_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIA_negPS10G_1_A_V_readaddr,
        doutb     => IL_L1PHIA_negPS10G_1_A_V_dout,
        sync_nent => IL_L1PHIA_negPS10G_1_A_start,
        nent_o    => IL_L1PHIA_negPS10G_1_A_AV_dout_nent
      );

    IL_L1PHIA_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIA_negPS10G_1_A_wea,
        addra     => IL_L1PHIA_negPS10G_1_A_writeaddr,
        dina      => IL_L1PHIA_negPS10G_1_A_din,
        wea_out       => IL_L1PHIA_negPS10G_1_A_wea_delay,
        addra_out     => IL_L1PHIA_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_L1PHIA_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIA_negPS10G_1_A_start
      );

    IL_L1PHIB_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIB_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIB_negPS10G_1_A_wea_delay,
        addra     => IL_L1PHIB_negPS10G_1_A_writeaddr_delay,
        dina      => IL_L1PHIB_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIB_negPS10G_1_A_V_readaddr,
        doutb     => IL_L1PHIB_negPS10G_1_A_V_dout,
        sync_nent => IL_L1PHIB_negPS10G_1_A_start,
        nent_o    => IL_L1PHIB_negPS10G_1_A_AV_dout_nent
      );

    IL_L1PHIB_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIB_negPS10G_1_A_wea,
        addra     => IL_L1PHIB_negPS10G_1_A_writeaddr,
        dina      => IL_L1PHIB_negPS10G_1_A_din,
        wea_out       => IL_L1PHIB_negPS10G_1_A_wea_delay,
        addra_out     => IL_L1PHIB_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_L1PHIB_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIB_negPS10G_1_A_start
      );

    IL_L1PHID_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHID_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHID_negPS10G_1_B_wea_delay,
        addra     => IL_L1PHID_negPS10G_1_B_writeaddr_delay,
        dina      => IL_L1PHID_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHID_negPS10G_1_B_V_readaddr,
        doutb     => IL_L1PHID_negPS10G_1_B_V_dout,
        sync_nent => IL_L1PHID_negPS10G_1_B_start,
        nent_o    => IL_L1PHID_negPS10G_1_B_AV_dout_nent
      );

    IL_L1PHID_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHID_negPS10G_1_B_wea,
        addra     => IL_L1PHID_negPS10G_1_B_writeaddr,
        dina      => IL_L1PHID_negPS10G_1_B_din,
        wea_out       => IL_L1PHID_negPS10G_1_B_wea_delay,
        addra_out     => IL_L1PHID_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_L1PHID_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHID_negPS10G_1_B_start
      );

    IL_L1PHIE_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIE_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIE_negPS10G_1_B_wea_delay,
        addra     => IL_L1PHIE_negPS10G_1_B_writeaddr_delay,
        dina      => IL_L1PHIE_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIE_negPS10G_1_B_V_readaddr,
        doutb     => IL_L1PHIE_negPS10G_1_B_V_dout,
        sync_nent => IL_L1PHIE_negPS10G_1_B_start,
        nent_o    => IL_L1PHIE_negPS10G_1_B_AV_dout_nent
      );

    IL_L1PHIE_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIE_negPS10G_1_B_wea,
        addra     => IL_L1PHIE_negPS10G_1_B_writeaddr,
        dina      => IL_L1PHIE_negPS10G_1_B_din,
        wea_out       => IL_L1PHIE_negPS10G_1_B_wea_delay,
        addra_out     => IL_L1PHIE_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_L1PHIE_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIE_negPS10G_1_B_start
      );

    IL_L1PHIF_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIF_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIF_negPS10G_1_B_wea_delay,
        addra     => IL_L1PHIF_negPS10G_1_B_writeaddr_delay,
        dina      => IL_L1PHIF_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIF_negPS10G_1_B_V_readaddr,
        doutb     => IL_L1PHIF_negPS10G_1_B_V_dout,
        sync_nent => IL_L1PHIF_negPS10G_1_B_start,
        nent_o    => IL_L1PHIF_negPS10G_1_B_AV_dout_nent
      );

    IL_L1PHIF_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIF_negPS10G_1_B_wea,
        addra     => IL_L1PHIF_negPS10G_1_B_writeaddr,
        dina      => IL_L1PHIF_negPS10G_1_B_din,
        wea_out       => IL_L1PHIF_negPS10G_1_B_wea_delay,
        addra_out     => IL_L1PHIF_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_L1PHIF_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIF_negPS10G_1_B_start
      );

    IL_L1PHIG_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIG_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIG_negPS10G_1_B_wea_delay,
        addra     => IL_L1PHIG_negPS10G_1_B_writeaddr_delay,
        dina      => IL_L1PHIG_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIG_negPS10G_1_B_V_readaddr,
        doutb     => IL_L1PHIG_negPS10G_1_B_V_dout,
        sync_nent => IL_L1PHIG_negPS10G_1_B_start,
        nent_o    => IL_L1PHIG_negPS10G_1_B_AV_dout_nent
      );

    IL_L1PHIG_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIG_negPS10G_1_B_wea,
        addra     => IL_L1PHIG_negPS10G_1_B_writeaddr,
        dina      => IL_L1PHIG_negPS10G_1_B_din,
        wea_out       => IL_L1PHIG_negPS10G_1_B_wea_delay,
        addra_out     => IL_L1PHIG_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_L1PHIG_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIG_negPS10G_1_B_start
      );

    IL_D1PHIA_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIA_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIA_negPS10G_1_A_wea_delay,
        addra     => IL_D1PHIA_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D1PHIA_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIA_negPS10G_1_A_V_readaddr,
        doutb     => IL_D1PHIA_negPS10G_1_A_V_dout,
        sync_nent => IL_D1PHIA_negPS10G_1_A_start,
        nent_o    => IL_D1PHIA_negPS10G_1_A_AV_dout_nent
      );

    IL_D1PHIA_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIA_negPS10G_1_A_wea,
        addra     => IL_D1PHIA_negPS10G_1_A_writeaddr,
        dina      => IL_D1PHIA_negPS10G_1_A_din,
        wea_out       => IL_D1PHIA_negPS10G_1_A_wea_delay,
        addra_out     => IL_D1PHIA_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D1PHIA_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIA_negPS10G_1_A_start
      );

    IL_D1PHIB_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_negPS10G_1_A_wea_delay,
        addra     => IL_D1PHIB_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D1PHIB_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_negPS10G_1_A_V_readaddr,
        doutb     => IL_D1PHIB_negPS10G_1_A_V_dout,
        sync_nent => IL_D1PHIB_negPS10G_1_A_start,
        nent_o    => IL_D1PHIB_negPS10G_1_A_AV_dout_nent
      );

    IL_D1PHIB_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_negPS10G_1_A_wea,
        addra     => IL_D1PHIB_negPS10G_1_A_writeaddr,
        dina      => IL_D1PHIB_negPS10G_1_A_din,
        wea_out       => IL_D1PHIB_negPS10G_1_A_wea_delay,
        addra_out     => IL_D1PHIB_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D1PHIB_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_negPS10G_1_A_start
      );

    IL_D1PHIB_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_negPS10G_1_B_wea_delay,
        addra     => IL_D1PHIB_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D1PHIB_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_negPS10G_1_B_V_readaddr,
        doutb     => IL_D1PHIB_negPS10G_1_B_V_dout,
        sync_nent => IL_D1PHIB_negPS10G_1_B_start,
        nent_o    => IL_D1PHIB_negPS10G_1_B_AV_dout_nent
      );

    IL_D1PHIB_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_negPS10G_1_B_wea,
        addra     => IL_D1PHIB_negPS10G_1_B_writeaddr,
        dina      => IL_D1PHIB_negPS10G_1_B_din,
        wea_out       => IL_D1PHIB_negPS10G_1_B_wea_delay,
        addra_out     => IL_D1PHIB_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D1PHIB_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_negPS10G_1_B_start
      );

    IL_D1PHIC_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_negPS10G_1_A_wea_delay,
        addra     => IL_D1PHIC_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D1PHIC_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_negPS10G_1_A_V_readaddr,
        doutb     => IL_D1PHIC_negPS10G_1_A_V_dout,
        sync_nent => IL_D1PHIC_negPS10G_1_A_start,
        nent_o    => IL_D1PHIC_negPS10G_1_A_AV_dout_nent
      );

    IL_D1PHIC_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_negPS10G_1_A_wea,
        addra     => IL_D1PHIC_negPS10G_1_A_writeaddr,
        dina      => IL_D1PHIC_negPS10G_1_A_din,
        wea_out       => IL_D1PHIC_negPS10G_1_A_wea_delay,
        addra_out     => IL_D1PHIC_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D1PHIC_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_negPS10G_1_A_start
      );

    IL_D1PHIC_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_negPS10G_1_B_wea_delay,
        addra     => IL_D1PHIC_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D1PHIC_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_negPS10G_1_B_V_readaddr,
        doutb     => IL_D1PHIC_negPS10G_1_B_V_dout,
        sync_nent => IL_D1PHIC_negPS10G_1_B_start,
        nent_o    => IL_D1PHIC_negPS10G_1_B_AV_dout_nent
      );

    IL_D1PHIC_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_negPS10G_1_B_wea,
        addra     => IL_D1PHIC_negPS10G_1_B_writeaddr,
        dina      => IL_D1PHIC_negPS10G_1_B_din,
        wea_out       => IL_D1PHIC_negPS10G_1_B_wea_delay,
        addra_out     => IL_D1PHIC_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D1PHIC_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_negPS10G_1_B_start
      );

    IL_D1PHID_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHID_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHID_negPS10G_1_B_wea_delay,
        addra     => IL_D1PHID_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D1PHID_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHID_negPS10G_1_B_V_readaddr,
        doutb     => IL_D1PHID_negPS10G_1_B_V_dout,
        sync_nent => IL_D1PHID_negPS10G_1_B_start,
        nent_o    => IL_D1PHID_negPS10G_1_B_AV_dout_nent
      );

    IL_D1PHID_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHID_negPS10G_1_B_wea,
        addra     => IL_D1PHID_negPS10G_1_B_writeaddr,
        dina      => IL_D1PHID_negPS10G_1_B_din,
        wea_out       => IL_D1PHID_negPS10G_1_B_wea_delay,
        addra_out     => IL_D1PHID_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D1PHID_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHID_negPS10G_1_B_start
      );

    IL_D3PHIA_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIA_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIA_negPS10G_1_A_wea_delay,
        addra     => IL_D3PHIA_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D3PHIA_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIA_negPS10G_1_A_V_readaddr,
        doutb     => IL_D3PHIA_negPS10G_1_A_V_dout,
        sync_nent => IL_D3PHIA_negPS10G_1_A_start,
        nent_o    => IL_D3PHIA_negPS10G_1_A_AV_dout_nent
      );

    IL_D3PHIA_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIA_negPS10G_1_A_wea,
        addra     => IL_D3PHIA_negPS10G_1_A_writeaddr,
        dina      => IL_D3PHIA_negPS10G_1_A_din,
        wea_out       => IL_D3PHIA_negPS10G_1_A_wea_delay,
        addra_out     => IL_D3PHIA_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D3PHIA_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIA_negPS10G_1_A_start
      );

    IL_D3PHIB_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_negPS10G_1_A_wea_delay,
        addra     => IL_D3PHIB_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D3PHIB_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_negPS10G_1_A_V_readaddr,
        doutb     => IL_D3PHIB_negPS10G_1_A_V_dout,
        sync_nent => IL_D3PHIB_negPS10G_1_A_start,
        nent_o    => IL_D3PHIB_negPS10G_1_A_AV_dout_nent
      );

    IL_D3PHIB_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_negPS10G_1_A_wea,
        addra     => IL_D3PHIB_negPS10G_1_A_writeaddr,
        dina      => IL_D3PHIB_negPS10G_1_A_din,
        wea_out       => IL_D3PHIB_negPS10G_1_A_wea_delay,
        addra_out     => IL_D3PHIB_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D3PHIB_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_negPS10G_1_A_start
      );

    IL_D3PHIB_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_negPS10G_1_B_wea_delay,
        addra     => IL_D3PHIB_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D3PHIB_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_negPS10G_1_B_V_readaddr,
        doutb     => IL_D3PHIB_negPS10G_1_B_V_dout,
        sync_nent => IL_D3PHIB_negPS10G_1_B_start,
        nent_o    => IL_D3PHIB_negPS10G_1_B_AV_dout_nent
      );

    IL_D3PHIB_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_negPS10G_1_B_wea,
        addra     => IL_D3PHIB_negPS10G_1_B_writeaddr,
        dina      => IL_D3PHIB_negPS10G_1_B_din,
        wea_out       => IL_D3PHIB_negPS10G_1_B_wea_delay,
        addra_out     => IL_D3PHIB_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D3PHIB_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_negPS10G_1_B_start
      );

    IL_D3PHIC_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_negPS10G_1_A_wea_delay,
        addra     => IL_D3PHIC_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D3PHIC_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_negPS10G_1_A_V_readaddr,
        doutb     => IL_D3PHIC_negPS10G_1_A_V_dout,
        sync_nent => IL_D3PHIC_negPS10G_1_A_start,
        nent_o    => IL_D3PHIC_negPS10G_1_A_AV_dout_nent
      );

    IL_D3PHIC_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_negPS10G_1_A_wea,
        addra     => IL_D3PHIC_negPS10G_1_A_writeaddr,
        dina      => IL_D3PHIC_negPS10G_1_A_din,
        wea_out       => IL_D3PHIC_negPS10G_1_A_wea_delay,
        addra_out     => IL_D3PHIC_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D3PHIC_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_negPS10G_1_A_start
      );

    IL_D3PHIC_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_negPS10G_1_B_wea_delay,
        addra     => IL_D3PHIC_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D3PHIC_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_negPS10G_1_B_V_readaddr,
        doutb     => IL_D3PHIC_negPS10G_1_B_V_dout,
        sync_nent => IL_D3PHIC_negPS10G_1_B_start,
        nent_o    => IL_D3PHIC_negPS10G_1_B_AV_dout_nent
      );

    IL_D3PHIC_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_negPS10G_1_B_wea,
        addra     => IL_D3PHIC_negPS10G_1_B_writeaddr,
        dina      => IL_D3PHIC_negPS10G_1_B_din,
        wea_out       => IL_D3PHIC_negPS10G_1_B_wea_delay,
        addra_out     => IL_D3PHIC_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D3PHIC_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_negPS10G_1_B_start
      );

    IL_D3PHID_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHID_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHID_negPS10G_1_B_wea_delay,
        addra     => IL_D3PHID_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D3PHID_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHID_negPS10G_1_B_V_readaddr,
        doutb     => IL_D3PHID_negPS10G_1_B_V_dout,
        sync_nent => IL_D3PHID_negPS10G_1_B_start,
        nent_o    => IL_D3PHID_negPS10G_1_B_AV_dout_nent
      );

    IL_D3PHID_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHID_negPS10G_1_B_wea,
        addra     => IL_D3PHID_negPS10G_1_B_writeaddr,
        dina      => IL_D3PHID_negPS10G_1_B_din,
        wea_out       => IL_D3PHID_negPS10G_1_B_wea_delay,
        addra_out     => IL_D3PHID_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D3PHID_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHID_negPS10G_1_B_start
      );

    IL_D5PHIA_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIA_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIA_negPS10G_1_A_wea_delay,
        addra     => IL_D5PHIA_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D5PHIA_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIA_negPS10G_1_A_V_readaddr,
        doutb     => IL_D5PHIA_negPS10G_1_A_V_dout,
        sync_nent => IL_D5PHIA_negPS10G_1_A_start,
        nent_o    => IL_D5PHIA_negPS10G_1_A_AV_dout_nent
      );

    IL_D5PHIA_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIA_negPS10G_1_A_wea,
        addra     => IL_D5PHIA_negPS10G_1_A_writeaddr,
        dina      => IL_D5PHIA_negPS10G_1_A_din,
        wea_out       => IL_D5PHIA_negPS10G_1_A_wea_delay,
        addra_out     => IL_D5PHIA_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D5PHIA_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIA_negPS10G_1_A_start
      );

    IL_D5PHIB_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_negPS10G_1_A_wea_delay,
        addra     => IL_D5PHIB_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D5PHIB_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_negPS10G_1_A_V_readaddr,
        doutb     => IL_D5PHIB_negPS10G_1_A_V_dout,
        sync_nent => IL_D5PHIB_negPS10G_1_A_start,
        nent_o    => IL_D5PHIB_negPS10G_1_A_AV_dout_nent
      );

    IL_D5PHIB_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_negPS10G_1_A_wea,
        addra     => IL_D5PHIB_negPS10G_1_A_writeaddr,
        dina      => IL_D5PHIB_negPS10G_1_A_din,
        wea_out       => IL_D5PHIB_negPS10G_1_A_wea_delay,
        addra_out     => IL_D5PHIB_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D5PHIB_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_negPS10G_1_A_start
      );

    IL_D5PHIB_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_negPS10G_1_B_wea_delay,
        addra     => IL_D5PHIB_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D5PHIB_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_negPS10G_1_B_V_readaddr,
        doutb     => IL_D5PHIB_negPS10G_1_B_V_dout,
        sync_nent => IL_D5PHIB_negPS10G_1_B_start,
        nent_o    => IL_D5PHIB_negPS10G_1_B_AV_dout_nent
      );

    IL_D5PHIB_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_negPS10G_1_B_wea,
        addra     => IL_D5PHIB_negPS10G_1_B_writeaddr,
        dina      => IL_D5PHIB_negPS10G_1_B_din,
        wea_out       => IL_D5PHIB_negPS10G_1_B_wea_delay,
        addra_out     => IL_D5PHIB_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D5PHIB_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_negPS10G_1_B_start
      );

    IL_D5PHIC_negPS10G_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_negPS10G_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_negPS10G_1_A_wea_delay,
        addra     => IL_D5PHIC_negPS10G_1_A_writeaddr_delay,
        dina      => IL_D5PHIC_negPS10G_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_negPS10G_1_A_V_readaddr,
        doutb     => IL_D5PHIC_negPS10G_1_A_V_dout,
        sync_nent => IL_D5PHIC_negPS10G_1_A_start,
        nent_o    => IL_D5PHIC_negPS10G_1_A_AV_dout_nent
      );

    IL_D5PHIC_negPS10G_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_negPS10G_1_A_wea,
        addra     => IL_D5PHIC_negPS10G_1_A_writeaddr,
        dina      => IL_D5PHIC_negPS10G_1_A_din,
        wea_out       => IL_D5PHIC_negPS10G_1_A_wea_delay,
        addra_out     => IL_D5PHIC_negPS10G_1_A_writeaddr_delay,
        dina_out      => IL_D5PHIC_negPS10G_1_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_negPS10G_1_A_start
      );

    IL_D5PHIC_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_negPS10G_1_B_wea_delay,
        addra     => IL_D5PHIC_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D5PHIC_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_negPS10G_1_B_V_readaddr,
        doutb     => IL_D5PHIC_negPS10G_1_B_V_dout,
        sync_nent => IL_D5PHIC_negPS10G_1_B_start,
        nent_o    => IL_D5PHIC_negPS10G_1_B_AV_dout_nent
      );

    IL_D5PHIC_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_negPS10G_1_B_wea,
        addra     => IL_D5PHIC_negPS10G_1_B_writeaddr,
        dina      => IL_D5PHIC_negPS10G_1_B_din,
        wea_out       => IL_D5PHIC_negPS10G_1_B_wea_delay,
        addra_out     => IL_D5PHIC_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D5PHIC_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_negPS10G_1_B_start
      );

    IL_D5PHID_negPS10G_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHID_negPS10G_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHID_negPS10G_1_B_wea_delay,
        addra     => IL_D5PHID_negPS10G_1_B_writeaddr_delay,
        dina      => IL_D5PHID_negPS10G_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHID_negPS10G_1_B_V_readaddr,
        doutb     => IL_D5PHID_negPS10G_1_B_V_dout,
        sync_nent => IL_D5PHID_negPS10G_1_B_start,
        nent_o    => IL_D5PHID_negPS10G_1_B_AV_dout_nent
      );

    IL_D5PHID_negPS10G_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHID_negPS10G_1_B_wea,
        addra     => IL_D5PHID_negPS10G_1_B_writeaddr,
        dina      => IL_D5PHID_negPS10G_1_B_din,
        wea_out       => IL_D5PHID_negPS10G_1_B_wea_delay,
        addra_out     => IL_D5PHID_negPS10G_1_B_writeaddr_delay,
        dina_out      => IL_D5PHID_negPS10G_1_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHID_negPS10G_1_B_start
      );

    IL_L1PHIA_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIA_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIA_negPS10G_2_A_wea_delay,
        addra     => IL_L1PHIA_negPS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIA_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIA_negPS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIA_negPS10G_2_A_V_dout,
        sync_nent => IL_L1PHIA_negPS10G_2_A_start,
        nent_o    => IL_L1PHIA_negPS10G_2_A_AV_dout_nent
      );

    IL_L1PHIA_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIA_negPS10G_2_A_wea,
        addra     => IL_L1PHIA_negPS10G_2_A_writeaddr,
        dina      => IL_L1PHIA_negPS10G_2_A_din,
        wea_out       => IL_L1PHIA_negPS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIA_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIA_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIA_negPS10G_2_A_start
      );

    IL_L1PHIB_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIB_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIB_negPS10G_2_A_wea_delay,
        addra     => IL_L1PHIB_negPS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIB_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIB_negPS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIB_negPS10G_2_A_V_dout,
        sync_nent => IL_L1PHIB_negPS10G_2_A_start,
        nent_o    => IL_L1PHIB_negPS10G_2_A_AV_dout_nent
      );

    IL_L1PHIB_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIB_negPS10G_2_A_wea,
        addra     => IL_L1PHIB_negPS10G_2_A_writeaddr,
        dina      => IL_L1PHIB_negPS10G_2_A_din,
        wea_out       => IL_L1PHIB_negPS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIB_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIB_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIB_negPS10G_2_A_start
      );

    IL_L1PHIC_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIC_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIC_negPS10G_2_A_wea_delay,
        addra     => IL_L1PHIC_negPS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIC_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIC_negPS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIC_negPS10G_2_A_V_dout,
        sync_nent => IL_L1PHIC_negPS10G_2_A_start,
        nent_o    => IL_L1PHIC_negPS10G_2_A_AV_dout_nent
      );

    IL_L1PHIC_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIC_negPS10G_2_A_wea,
        addra     => IL_L1PHIC_negPS10G_2_A_writeaddr,
        dina      => IL_L1PHIC_negPS10G_2_A_din,
        wea_out       => IL_L1PHIC_negPS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIC_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIC_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIC_negPS10G_2_A_start
      );

    IL_L1PHID_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHID_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHID_negPS10G_2_A_wea_delay,
        addra     => IL_L1PHID_negPS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHID_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHID_negPS10G_2_A_V_readaddr,
        doutb     => IL_L1PHID_negPS10G_2_A_V_dout,
        sync_nent => IL_L1PHID_negPS10G_2_A_start,
        nent_o    => IL_L1PHID_negPS10G_2_A_AV_dout_nent
      );

    IL_L1PHID_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHID_negPS10G_2_A_wea,
        addra     => IL_L1PHID_negPS10G_2_A_writeaddr,
        dina      => IL_L1PHID_negPS10G_2_A_din,
        wea_out       => IL_L1PHID_negPS10G_2_A_wea_delay,
        addra_out     => IL_L1PHID_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHID_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHID_negPS10G_2_A_start
      );

    IL_L1PHID_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHID_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHID_negPS10G_2_B_wea_delay,
        addra     => IL_L1PHID_negPS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHID_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHID_negPS10G_2_B_V_readaddr,
        doutb     => IL_L1PHID_negPS10G_2_B_V_dout,
        sync_nent => IL_L1PHID_negPS10G_2_B_start,
        nent_o    => IL_L1PHID_negPS10G_2_B_AV_dout_nent
      );

    IL_L1PHID_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHID_negPS10G_2_B_wea,
        addra     => IL_L1PHID_negPS10G_2_B_writeaddr,
        dina      => IL_L1PHID_negPS10G_2_B_din,
        wea_out       => IL_L1PHID_negPS10G_2_B_wea_delay,
        addra_out     => IL_L1PHID_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHID_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHID_negPS10G_2_B_start
      );

    IL_L1PHIE_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIE_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIE_negPS10G_2_A_wea_delay,
        addra     => IL_L1PHIE_negPS10G_2_A_writeaddr_delay,
        dina      => IL_L1PHIE_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIE_negPS10G_2_A_V_readaddr,
        doutb     => IL_L1PHIE_negPS10G_2_A_V_dout,
        sync_nent => IL_L1PHIE_negPS10G_2_A_start,
        nent_o    => IL_L1PHIE_negPS10G_2_A_AV_dout_nent
      );

    IL_L1PHIE_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIE_negPS10G_2_A_wea,
        addra     => IL_L1PHIE_negPS10G_2_A_writeaddr,
        dina      => IL_L1PHIE_negPS10G_2_A_din,
        wea_out       => IL_L1PHIE_negPS10G_2_A_wea_delay,
        addra_out     => IL_L1PHIE_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_L1PHIE_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_L1PHIE_negPS10G_2_A_start
      );

    IL_L1PHIE_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIE_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIE_negPS10G_2_B_wea_delay,
        addra     => IL_L1PHIE_negPS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIE_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIE_negPS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIE_negPS10G_2_B_V_dout,
        sync_nent => IL_L1PHIE_negPS10G_2_B_start,
        nent_o    => IL_L1PHIE_negPS10G_2_B_AV_dout_nent
      );

    IL_L1PHIE_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIE_negPS10G_2_B_wea,
        addra     => IL_L1PHIE_negPS10G_2_B_writeaddr,
        dina      => IL_L1PHIE_negPS10G_2_B_din,
        wea_out       => IL_L1PHIE_negPS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIE_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIE_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIE_negPS10G_2_B_start
      );

    IL_L1PHIF_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIF_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIF_negPS10G_2_B_wea_delay,
        addra     => IL_L1PHIF_negPS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIF_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIF_negPS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIF_negPS10G_2_B_V_dout,
        sync_nent => IL_L1PHIF_negPS10G_2_B_start,
        nent_o    => IL_L1PHIF_negPS10G_2_B_AV_dout_nent
      );

    IL_L1PHIF_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIF_negPS10G_2_B_wea,
        addra     => IL_L1PHIF_negPS10G_2_B_writeaddr,
        dina      => IL_L1PHIF_negPS10G_2_B_din,
        wea_out       => IL_L1PHIF_negPS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIF_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIF_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIF_negPS10G_2_B_start
      );

    IL_L1PHIG_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIG_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIG_negPS10G_2_B_wea_delay,
        addra     => IL_L1PHIG_negPS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIG_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIG_negPS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIG_negPS10G_2_B_V_dout,
        sync_nent => IL_L1PHIG_negPS10G_2_B_start,
        nent_o    => IL_L1PHIG_negPS10G_2_B_AV_dout_nent
      );

    IL_L1PHIG_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIG_negPS10G_2_B_wea,
        addra     => IL_L1PHIG_negPS10G_2_B_writeaddr,
        dina      => IL_L1PHIG_negPS10G_2_B_din,
        wea_out       => IL_L1PHIG_negPS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIG_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIG_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIG_negPS10G_2_B_start
      );

    IL_L1PHIH_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L1PHIH_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L1PHIH_negPS10G_2_B_wea_delay,
        addra     => IL_L1PHIH_negPS10G_2_B_writeaddr_delay,
        dina      => IL_L1PHIH_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L1PHIH_negPS10G_2_B_V_readaddr,
        doutb     => IL_L1PHIH_negPS10G_2_B_V_dout,
        sync_nent => IL_L1PHIH_negPS10G_2_B_start,
        nent_o    => IL_L1PHIH_negPS10G_2_B_AV_dout_nent
      );

    IL_L1PHIH_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L1PHIH_negPS10G_2_B_wea,
        addra     => IL_L1PHIH_negPS10G_2_B_writeaddr,
        dina      => IL_L1PHIH_negPS10G_2_B_din,
        wea_out       => IL_L1PHIH_negPS10G_2_B_wea_delay,
        addra_out     => IL_L1PHIH_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_L1PHIH_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_L1PHIH_negPS10G_2_B_start
      );

    IL_D2PHIA_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_negPS10G_2_A_wea_delay,
        addra     => IL_D2PHIA_negPS10G_2_A_writeaddr_delay,
        dina      => IL_D2PHIA_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_negPS10G_2_A_V_readaddr,
        doutb     => IL_D2PHIA_negPS10G_2_A_V_dout,
        sync_nent => IL_D2PHIA_negPS10G_2_A_start,
        nent_o    => IL_D2PHIA_negPS10G_2_A_AV_dout_nent
      );

    IL_D2PHIA_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_negPS10G_2_A_wea,
        addra     => IL_D2PHIA_negPS10G_2_A_writeaddr,
        dina      => IL_D2PHIA_negPS10G_2_A_din,
        wea_out       => IL_D2PHIA_negPS10G_2_A_wea_delay,
        addra_out     => IL_D2PHIA_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_negPS10G_2_A_start
      );

    IL_D2PHIB_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_negPS10G_2_A_wea_delay,
        addra     => IL_D2PHIB_negPS10G_2_A_writeaddr_delay,
        dina      => IL_D2PHIB_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_negPS10G_2_A_V_readaddr,
        doutb     => IL_D2PHIB_negPS10G_2_A_V_dout,
        sync_nent => IL_D2PHIB_negPS10G_2_A_start,
        nent_o    => IL_D2PHIB_negPS10G_2_A_AV_dout_nent
      );

    IL_D2PHIB_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_negPS10G_2_A_wea,
        addra     => IL_D2PHIB_negPS10G_2_A_writeaddr,
        dina      => IL_D2PHIB_negPS10G_2_A_din,
        wea_out       => IL_D2PHIB_negPS10G_2_A_wea_delay,
        addra_out     => IL_D2PHIB_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_negPS10G_2_A_start
      );

    IL_D2PHIB_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_negPS10G_2_B_wea_delay,
        addra     => IL_D2PHIB_negPS10G_2_B_writeaddr_delay,
        dina      => IL_D2PHIB_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_negPS10G_2_B_V_readaddr,
        doutb     => IL_D2PHIB_negPS10G_2_B_V_dout,
        sync_nent => IL_D2PHIB_negPS10G_2_B_start,
        nent_o    => IL_D2PHIB_negPS10G_2_B_AV_dout_nent
      );

    IL_D2PHIB_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_negPS10G_2_B_wea,
        addra     => IL_D2PHIB_negPS10G_2_B_writeaddr,
        dina      => IL_D2PHIB_negPS10G_2_B_din,
        wea_out       => IL_D2PHIB_negPS10G_2_B_wea_delay,
        addra_out     => IL_D2PHIB_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_negPS10G_2_B_start
      );

    IL_D2PHIC_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_negPS10G_2_A_wea_delay,
        addra     => IL_D2PHIC_negPS10G_2_A_writeaddr_delay,
        dina      => IL_D2PHIC_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_negPS10G_2_A_V_readaddr,
        doutb     => IL_D2PHIC_negPS10G_2_A_V_dout,
        sync_nent => IL_D2PHIC_negPS10G_2_A_start,
        nent_o    => IL_D2PHIC_negPS10G_2_A_AV_dout_nent
      );

    IL_D2PHIC_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_negPS10G_2_A_wea,
        addra     => IL_D2PHIC_negPS10G_2_A_writeaddr,
        dina      => IL_D2PHIC_negPS10G_2_A_din,
        wea_out       => IL_D2PHIC_negPS10G_2_A_wea_delay,
        addra_out     => IL_D2PHIC_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_negPS10G_2_A_start
      );

    IL_D2PHIC_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_negPS10G_2_B_wea_delay,
        addra     => IL_D2PHIC_negPS10G_2_B_writeaddr_delay,
        dina      => IL_D2PHIC_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_negPS10G_2_B_V_readaddr,
        doutb     => IL_D2PHIC_negPS10G_2_B_V_dout,
        sync_nent => IL_D2PHIC_negPS10G_2_B_start,
        nent_o    => IL_D2PHIC_negPS10G_2_B_AV_dout_nent
      );

    IL_D2PHIC_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_negPS10G_2_B_wea,
        addra     => IL_D2PHIC_negPS10G_2_B_writeaddr,
        dina      => IL_D2PHIC_negPS10G_2_B_din,
        wea_out       => IL_D2PHIC_negPS10G_2_B_wea_delay,
        addra_out     => IL_D2PHIC_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_negPS10G_2_B_start
      );

    IL_D2PHID_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_negPS10G_2_B_wea_delay,
        addra     => IL_D2PHID_negPS10G_2_B_writeaddr_delay,
        dina      => IL_D2PHID_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_negPS10G_2_B_V_readaddr,
        doutb     => IL_D2PHID_negPS10G_2_B_V_dout,
        sync_nent => IL_D2PHID_negPS10G_2_B_start,
        nent_o    => IL_D2PHID_negPS10G_2_B_AV_dout_nent
      );

    IL_D2PHID_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_negPS10G_2_B_wea,
        addra     => IL_D2PHID_negPS10G_2_B_writeaddr,
        dina      => IL_D2PHID_negPS10G_2_B_din,
        wea_out       => IL_D2PHID_negPS10G_2_B_wea_delay,
        addra_out     => IL_D2PHID_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_D2PHID_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_negPS10G_2_B_start
      );

    IL_D4PHIA_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIA_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIA_negPS10G_2_A_wea_delay,
        addra     => IL_D4PHIA_negPS10G_2_A_writeaddr_delay,
        dina      => IL_D4PHIA_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIA_negPS10G_2_A_V_readaddr,
        doutb     => IL_D4PHIA_negPS10G_2_A_V_dout,
        sync_nent => IL_D4PHIA_negPS10G_2_A_start,
        nent_o    => IL_D4PHIA_negPS10G_2_A_AV_dout_nent
      );

    IL_D4PHIA_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIA_negPS10G_2_A_wea,
        addra     => IL_D4PHIA_negPS10G_2_A_writeaddr,
        dina      => IL_D4PHIA_negPS10G_2_A_din,
        wea_out       => IL_D4PHIA_negPS10G_2_A_wea_delay,
        addra_out     => IL_D4PHIA_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIA_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIA_negPS10G_2_A_start
      );

    IL_D4PHIB_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_negPS10G_2_A_wea_delay,
        addra     => IL_D4PHIB_negPS10G_2_A_writeaddr_delay,
        dina      => IL_D4PHIB_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_negPS10G_2_A_V_readaddr,
        doutb     => IL_D4PHIB_negPS10G_2_A_V_dout,
        sync_nent => IL_D4PHIB_negPS10G_2_A_start,
        nent_o    => IL_D4PHIB_negPS10G_2_A_AV_dout_nent
      );

    IL_D4PHIB_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_negPS10G_2_A_wea,
        addra     => IL_D4PHIB_negPS10G_2_A_writeaddr,
        dina      => IL_D4PHIB_negPS10G_2_A_din,
        wea_out       => IL_D4PHIB_negPS10G_2_A_wea_delay,
        addra_out     => IL_D4PHIB_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIB_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_negPS10G_2_A_start
      );

    IL_D4PHIB_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_negPS10G_2_B_wea_delay,
        addra     => IL_D4PHIB_negPS10G_2_B_writeaddr_delay,
        dina      => IL_D4PHIB_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_negPS10G_2_B_V_readaddr,
        doutb     => IL_D4PHIB_negPS10G_2_B_V_dout,
        sync_nent => IL_D4PHIB_negPS10G_2_B_start,
        nent_o    => IL_D4PHIB_negPS10G_2_B_AV_dout_nent
      );

    IL_D4PHIB_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_negPS10G_2_B_wea,
        addra     => IL_D4PHIB_negPS10G_2_B_writeaddr,
        dina      => IL_D4PHIB_negPS10G_2_B_din,
        wea_out       => IL_D4PHIB_negPS10G_2_B_wea_delay,
        addra_out     => IL_D4PHIB_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIB_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_negPS10G_2_B_start
      );

    IL_D4PHIC_negPS10G_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_negPS10G_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_negPS10G_2_A_wea_delay,
        addra     => IL_D4PHIC_negPS10G_2_A_writeaddr_delay,
        dina      => IL_D4PHIC_negPS10G_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_negPS10G_2_A_V_readaddr,
        doutb     => IL_D4PHIC_negPS10G_2_A_V_dout,
        sync_nent => IL_D4PHIC_negPS10G_2_A_start,
        nent_o    => IL_D4PHIC_negPS10G_2_A_AV_dout_nent
      );

    IL_D4PHIC_negPS10G_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_negPS10G_2_A_wea,
        addra     => IL_D4PHIC_negPS10G_2_A_writeaddr,
        dina      => IL_D4PHIC_negPS10G_2_A_din,
        wea_out       => IL_D4PHIC_negPS10G_2_A_wea_delay,
        addra_out     => IL_D4PHIC_negPS10G_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIC_negPS10G_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_negPS10G_2_A_start
      );

    IL_D4PHIC_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_negPS10G_2_B_wea_delay,
        addra     => IL_D4PHIC_negPS10G_2_B_writeaddr_delay,
        dina      => IL_D4PHIC_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_negPS10G_2_B_V_readaddr,
        doutb     => IL_D4PHIC_negPS10G_2_B_V_dout,
        sync_nent => IL_D4PHIC_negPS10G_2_B_start,
        nent_o    => IL_D4PHIC_negPS10G_2_B_AV_dout_nent
      );

    IL_D4PHIC_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_negPS10G_2_B_wea,
        addra     => IL_D4PHIC_negPS10G_2_B_writeaddr,
        dina      => IL_D4PHIC_negPS10G_2_B_din,
        wea_out       => IL_D4PHIC_negPS10G_2_B_wea_delay,
        addra_out     => IL_D4PHIC_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIC_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_negPS10G_2_B_start
      );

    IL_D4PHID_negPS10G_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHID_negPS10G_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHID_negPS10G_2_B_wea_delay,
        addra     => IL_D4PHID_negPS10G_2_B_writeaddr_delay,
        dina      => IL_D4PHID_negPS10G_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHID_negPS10G_2_B_V_readaddr,
        doutb     => IL_D4PHID_negPS10G_2_B_V_dout,
        sync_nent => IL_D4PHID_negPS10G_2_B_start,
        nent_o    => IL_D4PHID_negPS10G_2_B_AV_dout_nent
      );

    IL_D4PHID_negPS10G_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHID_negPS10G_2_B_wea,
        addra     => IL_D4PHID_negPS10G_2_B_writeaddr,
        dina      => IL_D4PHID_negPS10G_2_B_din,
        wea_out       => IL_D4PHID_negPS10G_2_B_wea_delay,
        addra_out     => IL_D4PHID_negPS10G_2_B_writeaddr_delay,
        dina_out      => IL_D4PHID_negPS10G_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHID_negPS10G_2_B_start
      );

    IL_L2PHIA_negPS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIA_negPS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIA_negPS10G_3_A_wea_delay,
        addra     => IL_L2PHIA_negPS10G_3_A_writeaddr_delay,
        dina      => IL_L2PHIA_negPS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIA_negPS10G_3_A_V_readaddr,
        doutb     => IL_L2PHIA_negPS10G_3_A_V_dout,
        sync_nent => IL_L2PHIA_negPS10G_3_A_start,
        nent_o    => IL_L2PHIA_negPS10G_3_A_AV_dout_nent
      );

    IL_L2PHIA_negPS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIA_negPS10G_3_A_wea,
        addra     => IL_L2PHIA_negPS10G_3_A_writeaddr,
        dina      => IL_L2PHIA_negPS10G_3_A_din,
        wea_out       => IL_L2PHIA_negPS10G_3_A_wea_delay,
        addra_out     => IL_L2PHIA_negPS10G_3_A_writeaddr_delay,
        dina_out      => IL_L2PHIA_negPS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_L2PHIA_negPS10G_3_A_start
      );

    IL_L2PHIB_negPS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIB_negPS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIB_negPS10G_3_A_wea_delay,
        addra     => IL_L2PHIB_negPS10G_3_A_writeaddr_delay,
        dina      => IL_L2PHIB_negPS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIB_negPS10G_3_A_V_readaddr,
        doutb     => IL_L2PHIB_negPS10G_3_A_V_dout,
        sync_nent => IL_L2PHIB_negPS10G_3_A_start,
        nent_o    => IL_L2PHIB_negPS10G_3_A_AV_dout_nent
      );

    IL_L2PHIB_negPS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIB_negPS10G_3_A_wea,
        addra     => IL_L2PHIB_negPS10G_3_A_writeaddr,
        dina      => IL_L2PHIB_negPS10G_3_A_din,
        wea_out       => IL_L2PHIB_negPS10G_3_A_wea_delay,
        addra_out     => IL_L2PHIB_negPS10G_3_A_writeaddr_delay,
        dina_out      => IL_L2PHIB_negPS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_L2PHIB_negPS10G_3_A_start
      );

    IL_L2PHIB_negPS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIB_negPS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIB_negPS10G_3_B_wea_delay,
        addra     => IL_L2PHIB_negPS10G_3_B_writeaddr_delay,
        dina      => IL_L2PHIB_negPS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIB_negPS10G_3_B_V_readaddr,
        doutb     => IL_L2PHIB_negPS10G_3_B_V_dout,
        sync_nent => IL_L2PHIB_negPS10G_3_B_start,
        nent_o    => IL_L2PHIB_negPS10G_3_B_AV_dout_nent
      );

    IL_L2PHIB_negPS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIB_negPS10G_3_B_wea,
        addra     => IL_L2PHIB_negPS10G_3_B_writeaddr,
        dina      => IL_L2PHIB_negPS10G_3_B_din,
        wea_out       => IL_L2PHIB_negPS10G_3_B_wea_delay,
        addra_out     => IL_L2PHIB_negPS10G_3_B_writeaddr_delay,
        dina_out      => IL_L2PHIB_negPS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_L2PHIB_negPS10G_3_B_start
      );

    IL_L2PHIC_negPS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIC_negPS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIC_negPS10G_3_A_wea_delay,
        addra     => IL_L2PHIC_negPS10G_3_A_writeaddr_delay,
        dina      => IL_L2PHIC_negPS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIC_negPS10G_3_A_V_readaddr,
        doutb     => IL_L2PHIC_negPS10G_3_A_V_dout,
        sync_nent => IL_L2PHIC_negPS10G_3_A_start,
        nent_o    => IL_L2PHIC_negPS10G_3_A_AV_dout_nent
      );

    IL_L2PHIC_negPS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIC_negPS10G_3_A_wea,
        addra     => IL_L2PHIC_negPS10G_3_A_writeaddr,
        dina      => IL_L2PHIC_negPS10G_3_A_din,
        wea_out       => IL_L2PHIC_negPS10G_3_A_wea_delay,
        addra_out     => IL_L2PHIC_negPS10G_3_A_writeaddr_delay,
        dina_out      => IL_L2PHIC_negPS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_L2PHIC_negPS10G_3_A_start
      );

    IL_L2PHIC_negPS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHIC_negPS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHIC_negPS10G_3_B_wea_delay,
        addra     => IL_L2PHIC_negPS10G_3_B_writeaddr_delay,
        dina      => IL_L2PHIC_negPS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHIC_negPS10G_3_B_V_readaddr,
        doutb     => IL_L2PHIC_negPS10G_3_B_V_dout,
        sync_nent => IL_L2PHIC_negPS10G_3_B_start,
        nent_o    => IL_L2PHIC_negPS10G_3_B_AV_dout_nent
      );

    IL_L2PHIC_negPS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHIC_negPS10G_3_B_wea,
        addra     => IL_L2PHIC_negPS10G_3_B_writeaddr,
        dina      => IL_L2PHIC_negPS10G_3_B_din,
        wea_out       => IL_L2PHIC_negPS10G_3_B_wea_delay,
        addra_out     => IL_L2PHIC_negPS10G_3_B_writeaddr_delay,
        dina_out      => IL_L2PHIC_negPS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_L2PHIC_negPS10G_3_B_start
      );

    IL_L2PHID_negPS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L2PHID_negPS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L2PHID_negPS10G_3_B_wea_delay,
        addra     => IL_L2PHID_negPS10G_3_B_writeaddr_delay,
        dina      => IL_L2PHID_negPS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L2PHID_negPS10G_3_B_V_readaddr,
        doutb     => IL_L2PHID_negPS10G_3_B_V_dout,
        sync_nent => IL_L2PHID_negPS10G_3_B_start,
        nent_o    => IL_L2PHID_negPS10G_3_B_AV_dout_nent
      );

    IL_L2PHID_negPS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L2PHID_negPS10G_3_B_wea,
        addra     => IL_L2PHID_negPS10G_3_B_writeaddr,
        dina      => IL_L2PHID_negPS10G_3_B_din,
        wea_out       => IL_L2PHID_negPS10G_3_B_wea_delay,
        addra_out     => IL_L2PHID_negPS10G_3_B_writeaddr_delay,
        dina_out      => IL_L2PHID_negPS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_L2PHID_negPS10G_3_B_start
      );

    IL_D2PHIA_negPS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_negPS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_negPS10G_3_A_wea_delay,
        addra     => IL_D2PHIA_negPS10G_3_A_writeaddr_delay,
        dina      => IL_D2PHIA_negPS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_negPS10G_3_A_V_readaddr,
        doutb     => IL_D2PHIA_negPS10G_3_A_V_dout,
        sync_nent => IL_D2PHIA_negPS10G_3_A_start,
        nent_o    => IL_D2PHIA_negPS10G_3_A_AV_dout_nent
      );

    IL_D2PHIA_negPS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_negPS10G_3_A_wea,
        addra     => IL_D2PHIA_negPS10G_3_A_writeaddr,
        dina      => IL_D2PHIA_negPS10G_3_A_din,
        wea_out       => IL_D2PHIA_negPS10G_3_A_wea_delay,
        addra_out     => IL_D2PHIA_negPS10G_3_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_negPS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_negPS10G_3_A_start
      );

    IL_D2PHIB_negPS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_negPS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_negPS10G_3_A_wea_delay,
        addra     => IL_D2PHIB_negPS10G_3_A_writeaddr_delay,
        dina      => IL_D2PHIB_negPS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_negPS10G_3_A_V_readaddr,
        doutb     => IL_D2PHIB_negPS10G_3_A_V_dout,
        sync_nent => IL_D2PHIB_negPS10G_3_A_start,
        nent_o    => IL_D2PHIB_negPS10G_3_A_AV_dout_nent
      );

    IL_D2PHIB_negPS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_negPS10G_3_A_wea,
        addra     => IL_D2PHIB_negPS10G_3_A_writeaddr,
        dina      => IL_D2PHIB_negPS10G_3_A_din,
        wea_out       => IL_D2PHIB_negPS10G_3_A_wea_delay,
        addra_out     => IL_D2PHIB_negPS10G_3_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_negPS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_negPS10G_3_A_start
      );

    IL_D2PHIB_negPS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_negPS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_negPS10G_3_B_wea_delay,
        addra     => IL_D2PHIB_negPS10G_3_B_writeaddr_delay,
        dina      => IL_D2PHIB_negPS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_negPS10G_3_B_V_readaddr,
        doutb     => IL_D2PHIB_negPS10G_3_B_V_dout,
        sync_nent => IL_D2PHIB_negPS10G_3_B_start,
        nent_o    => IL_D2PHIB_negPS10G_3_B_AV_dout_nent
      );

    IL_D2PHIB_negPS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_negPS10G_3_B_wea,
        addra     => IL_D2PHIB_negPS10G_3_B_writeaddr,
        dina      => IL_D2PHIB_negPS10G_3_B_din,
        wea_out       => IL_D2PHIB_negPS10G_3_B_wea_delay,
        addra_out     => IL_D2PHIB_negPS10G_3_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_negPS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_negPS10G_3_B_start
      );

    IL_D2PHIC_negPS10G_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_negPS10G_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_negPS10G_3_A_wea_delay,
        addra     => IL_D2PHIC_negPS10G_3_A_writeaddr_delay,
        dina      => IL_D2PHIC_negPS10G_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_negPS10G_3_A_V_readaddr,
        doutb     => IL_D2PHIC_negPS10G_3_A_V_dout,
        sync_nent => IL_D2PHIC_negPS10G_3_A_start,
        nent_o    => IL_D2PHIC_negPS10G_3_A_AV_dout_nent
      );

    IL_D2PHIC_negPS10G_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_negPS10G_3_A_wea,
        addra     => IL_D2PHIC_negPS10G_3_A_writeaddr,
        dina      => IL_D2PHIC_negPS10G_3_A_din,
        wea_out       => IL_D2PHIC_negPS10G_3_A_wea_delay,
        addra_out     => IL_D2PHIC_negPS10G_3_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_negPS10G_3_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_negPS10G_3_A_start
      );

    IL_D2PHIC_negPS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_negPS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_negPS10G_3_B_wea_delay,
        addra     => IL_D2PHIC_negPS10G_3_B_writeaddr_delay,
        dina      => IL_D2PHIC_negPS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_negPS10G_3_B_V_readaddr,
        doutb     => IL_D2PHIC_negPS10G_3_B_V_dout,
        sync_nent => IL_D2PHIC_negPS10G_3_B_start,
        nent_o    => IL_D2PHIC_negPS10G_3_B_AV_dout_nent
      );

    IL_D2PHIC_negPS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_negPS10G_3_B_wea,
        addra     => IL_D2PHIC_negPS10G_3_B_writeaddr,
        dina      => IL_D2PHIC_negPS10G_3_B_din,
        wea_out       => IL_D2PHIC_negPS10G_3_B_wea_delay,
        addra_out     => IL_D2PHIC_negPS10G_3_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_negPS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_negPS10G_3_B_start
      );

    IL_D2PHID_negPS10G_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_negPS10G_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_negPS10G_3_B_wea_delay,
        addra     => IL_D2PHID_negPS10G_3_B_writeaddr_delay,
        dina      => IL_D2PHID_negPS10G_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_negPS10G_3_B_V_readaddr,
        doutb     => IL_D2PHID_negPS10G_3_B_V_dout,
        sync_nent => IL_D2PHID_negPS10G_3_B_start,
        nent_o    => IL_D2PHID_negPS10G_3_B_AV_dout_nent
      );

    IL_D2PHID_negPS10G_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_negPS10G_3_B_wea,
        addra     => IL_D2PHID_negPS10G_3_B_writeaddr,
        dina      => IL_D2PHID_negPS10G_3_B_din,
        wea_out       => IL_D2PHID_negPS10G_3_B_wea_delay,
        addra_out     => IL_D2PHID_negPS10G_3_B_writeaddr_delay,
        dina_out      => IL_D2PHID_negPS10G_3_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_negPS10G_3_B_start
      );

    IL_D1PHIA_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIA_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIA_negPS10G_4_A_wea_delay,
        addra     => IL_D1PHIA_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D1PHIA_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIA_negPS10G_4_A_V_readaddr,
        doutb     => IL_D1PHIA_negPS10G_4_A_V_dout,
        sync_nent => IL_D1PHIA_negPS10G_4_A_start,
        nent_o    => IL_D1PHIA_negPS10G_4_A_AV_dout_nent
      );

    IL_D1PHIA_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIA_negPS10G_4_A_wea,
        addra     => IL_D1PHIA_negPS10G_4_A_writeaddr,
        dina      => IL_D1PHIA_negPS10G_4_A_din,
        wea_out       => IL_D1PHIA_negPS10G_4_A_wea_delay,
        addra_out     => IL_D1PHIA_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D1PHIA_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIA_negPS10G_4_A_start
      );

    IL_D1PHIB_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_negPS10G_4_A_wea_delay,
        addra     => IL_D1PHIB_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D1PHIB_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_negPS10G_4_A_V_readaddr,
        doutb     => IL_D1PHIB_negPS10G_4_A_V_dout,
        sync_nent => IL_D1PHIB_negPS10G_4_A_start,
        nent_o    => IL_D1PHIB_negPS10G_4_A_AV_dout_nent
      );

    IL_D1PHIB_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_negPS10G_4_A_wea,
        addra     => IL_D1PHIB_negPS10G_4_A_writeaddr,
        dina      => IL_D1PHIB_negPS10G_4_A_din,
        wea_out       => IL_D1PHIB_negPS10G_4_A_wea_delay,
        addra_out     => IL_D1PHIB_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D1PHIB_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_negPS10G_4_A_start
      );

    IL_D1PHIB_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_negPS10G_4_B_wea_delay,
        addra     => IL_D1PHIB_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D1PHIB_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_negPS10G_4_B_V_readaddr,
        doutb     => IL_D1PHIB_negPS10G_4_B_V_dout,
        sync_nent => IL_D1PHIB_negPS10G_4_B_start,
        nent_o    => IL_D1PHIB_negPS10G_4_B_AV_dout_nent
      );

    IL_D1PHIB_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_negPS10G_4_B_wea,
        addra     => IL_D1PHIB_negPS10G_4_B_writeaddr,
        dina      => IL_D1PHIB_negPS10G_4_B_din,
        wea_out       => IL_D1PHIB_negPS10G_4_B_wea_delay,
        addra_out     => IL_D1PHIB_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D1PHIB_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_negPS10G_4_B_start
      );

    IL_D1PHIC_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_negPS10G_4_A_wea_delay,
        addra     => IL_D1PHIC_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D1PHIC_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_negPS10G_4_A_V_readaddr,
        doutb     => IL_D1PHIC_negPS10G_4_A_V_dout,
        sync_nent => IL_D1PHIC_negPS10G_4_A_start,
        nent_o    => IL_D1PHIC_negPS10G_4_A_AV_dout_nent
      );

    IL_D1PHIC_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_negPS10G_4_A_wea,
        addra     => IL_D1PHIC_negPS10G_4_A_writeaddr,
        dina      => IL_D1PHIC_negPS10G_4_A_din,
        wea_out       => IL_D1PHIC_negPS10G_4_A_wea_delay,
        addra_out     => IL_D1PHIC_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D1PHIC_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_negPS10G_4_A_start
      );

    IL_D1PHIC_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_negPS10G_4_B_wea_delay,
        addra     => IL_D1PHIC_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D1PHIC_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_negPS10G_4_B_V_readaddr,
        doutb     => IL_D1PHIC_negPS10G_4_B_V_dout,
        sync_nent => IL_D1PHIC_negPS10G_4_B_start,
        nent_o    => IL_D1PHIC_negPS10G_4_B_AV_dout_nent
      );

    IL_D1PHIC_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_negPS10G_4_B_wea,
        addra     => IL_D1PHIC_negPS10G_4_B_writeaddr,
        dina      => IL_D1PHIC_negPS10G_4_B_din,
        wea_out       => IL_D1PHIC_negPS10G_4_B_wea_delay,
        addra_out     => IL_D1PHIC_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D1PHIC_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_negPS10G_4_B_start
      );

    IL_D1PHID_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHID_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHID_negPS10G_4_B_wea_delay,
        addra     => IL_D1PHID_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D1PHID_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHID_negPS10G_4_B_V_readaddr,
        doutb     => IL_D1PHID_negPS10G_4_B_V_dout,
        sync_nent => IL_D1PHID_negPS10G_4_B_start,
        nent_o    => IL_D1PHID_negPS10G_4_B_AV_dout_nent
      );

    IL_D1PHID_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHID_negPS10G_4_B_wea,
        addra     => IL_D1PHID_negPS10G_4_B_writeaddr,
        dina      => IL_D1PHID_negPS10G_4_B_din,
        wea_out       => IL_D1PHID_negPS10G_4_B_wea_delay,
        addra_out     => IL_D1PHID_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D1PHID_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHID_negPS10G_4_B_start
      );

    IL_D3PHIA_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIA_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIA_negPS10G_4_A_wea_delay,
        addra     => IL_D3PHIA_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D3PHIA_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIA_negPS10G_4_A_V_readaddr,
        doutb     => IL_D3PHIA_negPS10G_4_A_V_dout,
        sync_nent => IL_D3PHIA_negPS10G_4_A_start,
        nent_o    => IL_D3PHIA_negPS10G_4_A_AV_dout_nent
      );

    IL_D3PHIA_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIA_negPS10G_4_A_wea,
        addra     => IL_D3PHIA_negPS10G_4_A_writeaddr,
        dina      => IL_D3PHIA_negPS10G_4_A_din,
        wea_out       => IL_D3PHIA_negPS10G_4_A_wea_delay,
        addra_out     => IL_D3PHIA_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIA_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIA_negPS10G_4_A_start
      );

    IL_D3PHIB_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_negPS10G_4_A_wea_delay,
        addra     => IL_D3PHIB_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D3PHIB_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_negPS10G_4_A_V_readaddr,
        doutb     => IL_D3PHIB_negPS10G_4_A_V_dout,
        sync_nent => IL_D3PHIB_negPS10G_4_A_start,
        nent_o    => IL_D3PHIB_negPS10G_4_A_AV_dout_nent
      );

    IL_D3PHIB_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_negPS10G_4_A_wea,
        addra     => IL_D3PHIB_negPS10G_4_A_writeaddr,
        dina      => IL_D3PHIB_negPS10G_4_A_din,
        wea_out       => IL_D3PHIB_negPS10G_4_A_wea_delay,
        addra_out     => IL_D3PHIB_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIB_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_negPS10G_4_A_start
      );

    IL_D3PHIB_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_negPS10G_4_B_wea_delay,
        addra     => IL_D3PHIB_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D3PHIB_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_negPS10G_4_B_V_readaddr,
        doutb     => IL_D3PHIB_negPS10G_4_B_V_dout,
        sync_nent => IL_D3PHIB_negPS10G_4_B_start,
        nent_o    => IL_D3PHIB_negPS10G_4_B_AV_dout_nent
      );

    IL_D3PHIB_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_negPS10G_4_B_wea,
        addra     => IL_D3PHIB_negPS10G_4_B_writeaddr,
        dina      => IL_D3PHIB_negPS10G_4_B_din,
        wea_out       => IL_D3PHIB_negPS10G_4_B_wea_delay,
        addra_out     => IL_D3PHIB_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIB_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_negPS10G_4_B_start
      );

    IL_D3PHIC_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_negPS10G_4_A_wea_delay,
        addra     => IL_D3PHIC_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D3PHIC_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_negPS10G_4_A_V_readaddr,
        doutb     => IL_D3PHIC_negPS10G_4_A_V_dout,
        sync_nent => IL_D3PHIC_negPS10G_4_A_start,
        nent_o    => IL_D3PHIC_negPS10G_4_A_AV_dout_nent
      );

    IL_D3PHIC_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_negPS10G_4_A_wea,
        addra     => IL_D3PHIC_negPS10G_4_A_writeaddr,
        dina      => IL_D3PHIC_negPS10G_4_A_din,
        wea_out       => IL_D3PHIC_negPS10G_4_A_wea_delay,
        addra_out     => IL_D3PHIC_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIC_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_negPS10G_4_A_start
      );

    IL_D3PHIC_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_negPS10G_4_B_wea_delay,
        addra     => IL_D3PHIC_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D3PHIC_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_negPS10G_4_B_V_readaddr,
        doutb     => IL_D3PHIC_negPS10G_4_B_V_dout,
        sync_nent => IL_D3PHIC_negPS10G_4_B_start,
        nent_o    => IL_D3PHIC_negPS10G_4_B_AV_dout_nent
      );

    IL_D3PHIC_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_negPS10G_4_B_wea,
        addra     => IL_D3PHIC_negPS10G_4_B_writeaddr,
        dina      => IL_D3PHIC_negPS10G_4_B_din,
        wea_out       => IL_D3PHIC_negPS10G_4_B_wea_delay,
        addra_out     => IL_D3PHIC_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIC_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_negPS10G_4_B_start
      );

    IL_D3PHID_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHID_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHID_negPS10G_4_B_wea_delay,
        addra     => IL_D3PHID_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D3PHID_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHID_negPS10G_4_B_V_readaddr,
        doutb     => IL_D3PHID_negPS10G_4_B_V_dout,
        sync_nent => IL_D3PHID_negPS10G_4_B_start,
        nent_o    => IL_D3PHID_negPS10G_4_B_AV_dout_nent
      );

    IL_D3PHID_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHID_negPS10G_4_B_wea,
        addra     => IL_D3PHID_negPS10G_4_B_writeaddr,
        dina      => IL_D3PHID_negPS10G_4_B_din,
        wea_out       => IL_D3PHID_negPS10G_4_B_wea_delay,
        addra_out     => IL_D3PHID_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D3PHID_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHID_negPS10G_4_B_start
      );

    IL_D5PHIA_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIA_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIA_negPS10G_4_A_wea_delay,
        addra     => IL_D5PHIA_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D5PHIA_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIA_negPS10G_4_A_V_readaddr,
        doutb     => IL_D5PHIA_negPS10G_4_A_V_dout,
        sync_nent => IL_D5PHIA_negPS10G_4_A_start,
        nent_o    => IL_D5PHIA_negPS10G_4_A_AV_dout_nent
      );

    IL_D5PHIA_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIA_negPS10G_4_A_wea,
        addra     => IL_D5PHIA_negPS10G_4_A_writeaddr,
        dina      => IL_D5PHIA_negPS10G_4_A_din,
        wea_out       => IL_D5PHIA_negPS10G_4_A_wea_delay,
        addra_out     => IL_D5PHIA_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D5PHIA_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIA_negPS10G_4_A_start
      );

    IL_D5PHIB_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_negPS10G_4_A_wea_delay,
        addra     => IL_D5PHIB_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D5PHIB_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_negPS10G_4_A_V_readaddr,
        doutb     => IL_D5PHIB_negPS10G_4_A_V_dout,
        sync_nent => IL_D5PHIB_negPS10G_4_A_start,
        nent_o    => IL_D5PHIB_negPS10G_4_A_AV_dout_nent
      );

    IL_D5PHIB_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_negPS10G_4_A_wea,
        addra     => IL_D5PHIB_negPS10G_4_A_writeaddr,
        dina      => IL_D5PHIB_negPS10G_4_A_din,
        wea_out       => IL_D5PHIB_negPS10G_4_A_wea_delay,
        addra_out     => IL_D5PHIB_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D5PHIB_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_negPS10G_4_A_start
      );

    IL_D5PHIB_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_negPS10G_4_B_wea_delay,
        addra     => IL_D5PHIB_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D5PHIB_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_negPS10G_4_B_V_readaddr,
        doutb     => IL_D5PHIB_negPS10G_4_B_V_dout,
        sync_nent => IL_D5PHIB_negPS10G_4_B_start,
        nent_o    => IL_D5PHIB_negPS10G_4_B_AV_dout_nent
      );

    IL_D5PHIB_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_negPS10G_4_B_wea,
        addra     => IL_D5PHIB_negPS10G_4_B_writeaddr,
        dina      => IL_D5PHIB_negPS10G_4_B_din,
        wea_out       => IL_D5PHIB_negPS10G_4_B_wea_delay,
        addra_out     => IL_D5PHIB_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D5PHIB_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_negPS10G_4_B_start
      );

    IL_D5PHIC_negPS10G_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_negPS10G_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_negPS10G_4_A_wea_delay,
        addra     => IL_D5PHIC_negPS10G_4_A_writeaddr_delay,
        dina      => IL_D5PHIC_negPS10G_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_negPS10G_4_A_V_readaddr,
        doutb     => IL_D5PHIC_negPS10G_4_A_V_dout,
        sync_nent => IL_D5PHIC_negPS10G_4_A_start,
        nent_o    => IL_D5PHIC_negPS10G_4_A_AV_dout_nent
      );

    IL_D5PHIC_negPS10G_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_negPS10G_4_A_wea,
        addra     => IL_D5PHIC_negPS10G_4_A_writeaddr,
        dina      => IL_D5PHIC_negPS10G_4_A_din,
        wea_out       => IL_D5PHIC_negPS10G_4_A_wea_delay,
        addra_out     => IL_D5PHIC_negPS10G_4_A_writeaddr_delay,
        dina_out      => IL_D5PHIC_negPS10G_4_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_negPS10G_4_A_start
      );

    IL_D5PHIC_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_negPS10G_4_B_wea_delay,
        addra     => IL_D5PHIC_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D5PHIC_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_negPS10G_4_B_V_readaddr,
        doutb     => IL_D5PHIC_negPS10G_4_B_V_dout,
        sync_nent => IL_D5PHIC_negPS10G_4_B_start,
        nent_o    => IL_D5PHIC_negPS10G_4_B_AV_dout_nent
      );

    IL_D5PHIC_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_negPS10G_4_B_wea,
        addra     => IL_D5PHIC_negPS10G_4_B_writeaddr,
        dina      => IL_D5PHIC_negPS10G_4_B_din,
        wea_out       => IL_D5PHIC_negPS10G_4_B_wea_delay,
        addra_out     => IL_D5PHIC_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D5PHIC_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_negPS10G_4_B_start
      );

    IL_D5PHID_negPS10G_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHID_negPS10G_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHID_negPS10G_4_B_wea_delay,
        addra     => IL_D5PHID_negPS10G_4_B_writeaddr_delay,
        dina      => IL_D5PHID_negPS10G_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHID_negPS10G_4_B_V_readaddr,
        doutb     => IL_D5PHID_negPS10G_4_B_V_dout,
        sync_nent => IL_D5PHID_negPS10G_4_B_start,
        nent_o    => IL_D5PHID_negPS10G_4_B_AV_dout_nent
      );

    IL_D5PHID_negPS10G_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHID_negPS10G_4_B_wea,
        addra     => IL_D5PHID_negPS10G_4_B_writeaddr,
        dina      => IL_D5PHID_negPS10G_4_B_din,
        wea_out       => IL_D5PHID_negPS10G_4_B_wea_delay,
        addra_out     => IL_D5PHID_negPS10G_4_B_writeaddr_delay,
        dina_out      => IL_D5PHID_negPS10G_4_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHID_negPS10G_4_B_start
      );

    IL_L3PHIA_negPS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIA_negPS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIA_negPS_1_A_wea_delay,
        addra     => IL_L3PHIA_negPS_1_A_writeaddr_delay,
        dina      => IL_L3PHIA_negPS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIA_negPS_1_A_V_readaddr,
        doutb     => IL_L3PHIA_negPS_1_A_V_dout,
        sync_nent => IL_L3PHIA_negPS_1_A_start,
        nent_o    => IL_L3PHIA_negPS_1_A_AV_dout_nent
      );

    IL_L3PHIA_negPS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIA_negPS_1_A_wea,
        addra     => IL_L3PHIA_negPS_1_A_writeaddr,
        dina      => IL_L3PHIA_negPS_1_A_din,
        wea_out       => IL_L3PHIA_negPS_1_A_wea_delay,
        addra_out     => IL_L3PHIA_negPS_1_A_writeaddr_delay,
        dina_out      => IL_L3PHIA_negPS_1_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIA_negPS_1_A_start
      );

    IL_L3PHIB_negPS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIB_negPS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIB_negPS_1_A_wea_delay,
        addra     => IL_L3PHIB_negPS_1_A_writeaddr_delay,
        dina      => IL_L3PHIB_negPS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIB_negPS_1_A_V_readaddr,
        doutb     => IL_L3PHIB_negPS_1_A_V_dout,
        sync_nent => IL_L3PHIB_negPS_1_A_start,
        nent_o    => IL_L3PHIB_negPS_1_A_AV_dout_nent
      );

    IL_L3PHIB_negPS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIB_negPS_1_A_wea,
        addra     => IL_L3PHIB_negPS_1_A_writeaddr,
        dina      => IL_L3PHIB_negPS_1_A_din,
        wea_out       => IL_L3PHIB_negPS_1_A_wea_delay,
        addra_out     => IL_L3PHIB_negPS_1_A_writeaddr_delay,
        dina_out      => IL_L3PHIB_negPS_1_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIB_negPS_1_A_start
      );

    IL_L3PHIB_negPS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIB_negPS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIB_negPS_1_B_wea_delay,
        addra     => IL_L3PHIB_negPS_1_B_writeaddr_delay,
        dina      => IL_L3PHIB_negPS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIB_negPS_1_B_V_readaddr,
        doutb     => IL_L3PHIB_negPS_1_B_V_dout,
        sync_nent => IL_L3PHIB_negPS_1_B_start,
        nent_o    => IL_L3PHIB_negPS_1_B_AV_dout_nent
      );

    IL_L3PHIB_negPS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIB_negPS_1_B_wea,
        addra     => IL_L3PHIB_negPS_1_B_writeaddr,
        dina      => IL_L3PHIB_negPS_1_B_din,
        wea_out       => IL_L3PHIB_negPS_1_B_wea_delay,
        addra_out     => IL_L3PHIB_negPS_1_B_writeaddr_delay,
        dina_out      => IL_L3PHIB_negPS_1_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHIB_negPS_1_B_start
      );

    IL_L3PHIC_negPS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIC_negPS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIC_negPS_1_B_wea_delay,
        addra     => IL_L3PHIC_negPS_1_B_writeaddr_delay,
        dina      => IL_L3PHIC_negPS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIC_negPS_1_B_V_readaddr,
        doutb     => IL_L3PHIC_negPS_1_B_V_dout,
        sync_nent => IL_L3PHIC_negPS_1_B_start,
        nent_o    => IL_L3PHIC_negPS_1_B_AV_dout_nent
      );

    IL_L3PHIC_negPS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIC_negPS_1_B_wea,
        addra     => IL_L3PHIC_negPS_1_B_writeaddr,
        dina      => IL_L3PHIC_negPS_1_B_din,
        wea_out       => IL_L3PHIC_negPS_1_B_wea_delay,
        addra_out     => IL_L3PHIC_negPS_1_B_writeaddr_delay,
        dina_out      => IL_L3PHIC_negPS_1_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHIC_negPS_1_B_start
      );

    IL_L3PHID_negPS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHID_negPS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHID_negPS_1_B_wea_delay,
        addra     => IL_L3PHID_negPS_1_B_writeaddr_delay,
        dina      => IL_L3PHID_negPS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHID_negPS_1_B_V_readaddr,
        doutb     => IL_L3PHID_negPS_1_B_V_dout,
        sync_nent => IL_L3PHID_negPS_1_B_start,
        nent_o    => IL_L3PHID_negPS_1_B_AV_dout_nent
      );

    IL_L3PHID_negPS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHID_negPS_1_B_wea,
        addra     => IL_L3PHID_negPS_1_B_writeaddr,
        dina      => IL_L3PHID_negPS_1_B_din,
        wea_out       => IL_L3PHID_negPS_1_B_wea_delay,
        addra_out     => IL_L3PHID_negPS_1_B_writeaddr_delay,
        dina_out      => IL_L3PHID_negPS_1_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHID_negPS_1_B_start
      );

    IL_D2PHIA_negPS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_negPS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_negPS_1_A_wea_delay,
        addra     => IL_D2PHIA_negPS_1_A_writeaddr_delay,
        dina      => IL_D2PHIA_negPS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_negPS_1_A_V_readaddr,
        doutb     => IL_D2PHIA_negPS_1_A_V_dout,
        sync_nent => IL_D2PHIA_negPS_1_A_start,
        nent_o    => IL_D2PHIA_negPS_1_A_AV_dout_nent
      );

    IL_D2PHIA_negPS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_negPS_1_A_wea,
        addra     => IL_D2PHIA_negPS_1_A_writeaddr,
        dina      => IL_D2PHIA_negPS_1_A_din,
        wea_out       => IL_D2PHIA_negPS_1_A_wea_delay,
        addra_out     => IL_D2PHIA_negPS_1_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_negPS_1_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_negPS_1_A_start
      );

    IL_D2PHIB_negPS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_negPS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_negPS_1_A_wea_delay,
        addra     => IL_D2PHIB_negPS_1_A_writeaddr_delay,
        dina      => IL_D2PHIB_negPS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_negPS_1_A_V_readaddr,
        doutb     => IL_D2PHIB_negPS_1_A_V_dout,
        sync_nent => IL_D2PHIB_negPS_1_A_start,
        nent_o    => IL_D2PHIB_negPS_1_A_AV_dout_nent
      );

    IL_D2PHIB_negPS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_negPS_1_A_wea,
        addra     => IL_D2PHIB_negPS_1_A_writeaddr,
        dina      => IL_D2PHIB_negPS_1_A_din,
        wea_out       => IL_D2PHIB_negPS_1_A_wea_delay,
        addra_out     => IL_D2PHIB_negPS_1_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_negPS_1_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_negPS_1_A_start
      );

    IL_D2PHIB_negPS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_negPS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_negPS_1_B_wea_delay,
        addra     => IL_D2PHIB_negPS_1_B_writeaddr_delay,
        dina      => IL_D2PHIB_negPS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_negPS_1_B_V_readaddr,
        doutb     => IL_D2PHIB_negPS_1_B_V_dout,
        sync_nent => IL_D2PHIB_negPS_1_B_start,
        nent_o    => IL_D2PHIB_negPS_1_B_AV_dout_nent
      );

    IL_D2PHIB_negPS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_negPS_1_B_wea,
        addra     => IL_D2PHIB_negPS_1_B_writeaddr,
        dina      => IL_D2PHIB_negPS_1_B_din,
        wea_out       => IL_D2PHIB_negPS_1_B_wea_delay,
        addra_out     => IL_D2PHIB_negPS_1_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_negPS_1_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_negPS_1_B_start
      );

    IL_D2PHIC_negPS_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_negPS_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_negPS_1_A_wea_delay,
        addra     => IL_D2PHIC_negPS_1_A_writeaddr_delay,
        dina      => IL_D2PHIC_negPS_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_negPS_1_A_V_readaddr,
        doutb     => IL_D2PHIC_negPS_1_A_V_dout,
        sync_nent => IL_D2PHIC_negPS_1_A_start,
        nent_o    => IL_D2PHIC_negPS_1_A_AV_dout_nent
      );

    IL_D2PHIC_negPS_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_negPS_1_A_wea,
        addra     => IL_D2PHIC_negPS_1_A_writeaddr,
        dina      => IL_D2PHIC_negPS_1_A_din,
        wea_out       => IL_D2PHIC_negPS_1_A_wea_delay,
        addra_out     => IL_D2PHIC_negPS_1_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_negPS_1_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_negPS_1_A_start
      );

    IL_D2PHIC_negPS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_negPS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_negPS_1_B_wea_delay,
        addra     => IL_D2PHIC_negPS_1_B_writeaddr_delay,
        dina      => IL_D2PHIC_negPS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_negPS_1_B_V_readaddr,
        doutb     => IL_D2PHIC_negPS_1_B_V_dout,
        sync_nent => IL_D2PHIC_negPS_1_B_start,
        nent_o    => IL_D2PHIC_negPS_1_B_AV_dout_nent
      );

    IL_D2PHIC_negPS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_negPS_1_B_wea,
        addra     => IL_D2PHIC_negPS_1_B_writeaddr,
        dina      => IL_D2PHIC_negPS_1_B_din,
        wea_out       => IL_D2PHIC_negPS_1_B_wea_delay,
        addra_out     => IL_D2PHIC_negPS_1_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_negPS_1_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_negPS_1_B_start
      );

    IL_D2PHID_negPS_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_negPS_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_negPS_1_B_wea_delay,
        addra     => IL_D2PHID_negPS_1_B_writeaddr_delay,
        dina      => IL_D2PHID_negPS_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_negPS_1_B_V_readaddr,
        doutb     => IL_D2PHID_negPS_1_B_V_dout,
        sync_nent => IL_D2PHID_negPS_1_B_start,
        nent_o    => IL_D2PHID_negPS_1_B_AV_dout_nent
      );

    IL_D2PHID_negPS_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_negPS_1_B_wea,
        addra     => IL_D2PHID_negPS_1_B_writeaddr,
        dina      => IL_D2PHID_negPS_1_B_din,
        wea_out       => IL_D2PHID_negPS_1_B_wea_delay,
        addra_out     => IL_D2PHID_negPS_1_B_writeaddr_delay,
        dina_out      => IL_D2PHID_negPS_1_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_negPS_1_B_start
      );

    IL_L3PHIA_negPS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIA_negPS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIA_negPS_2_A_wea_delay,
        addra     => IL_L3PHIA_negPS_2_A_writeaddr_delay,
        dina      => IL_L3PHIA_negPS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIA_negPS_2_A_V_readaddr,
        doutb     => IL_L3PHIA_negPS_2_A_V_dout,
        sync_nent => IL_L3PHIA_negPS_2_A_start,
        nent_o    => IL_L3PHIA_negPS_2_A_AV_dout_nent
      );

    IL_L3PHIA_negPS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIA_negPS_2_A_wea,
        addra     => IL_L3PHIA_negPS_2_A_writeaddr,
        dina      => IL_L3PHIA_negPS_2_A_din,
        wea_out       => IL_L3PHIA_negPS_2_A_wea_delay,
        addra_out     => IL_L3PHIA_negPS_2_A_writeaddr_delay,
        dina_out      => IL_L3PHIA_negPS_2_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIA_negPS_2_A_start
      );

    IL_L3PHIB_negPS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIB_negPS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIB_negPS_2_A_wea_delay,
        addra     => IL_L3PHIB_negPS_2_A_writeaddr_delay,
        dina      => IL_L3PHIB_negPS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIB_negPS_2_A_V_readaddr,
        doutb     => IL_L3PHIB_negPS_2_A_V_dout,
        sync_nent => IL_L3PHIB_negPS_2_A_start,
        nent_o    => IL_L3PHIB_negPS_2_A_AV_dout_nent
      );

    IL_L3PHIB_negPS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIB_negPS_2_A_wea,
        addra     => IL_L3PHIB_negPS_2_A_writeaddr,
        dina      => IL_L3PHIB_negPS_2_A_din,
        wea_out       => IL_L3PHIB_negPS_2_A_wea_delay,
        addra_out     => IL_L3PHIB_negPS_2_A_writeaddr_delay,
        dina_out      => IL_L3PHIB_negPS_2_A_din_delay,
        done       => IR_done,
        start      => IL_L3PHIB_negPS_2_A_start
      );

    IL_L3PHIB_negPS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIB_negPS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIB_negPS_2_B_wea_delay,
        addra     => IL_L3PHIB_negPS_2_B_writeaddr_delay,
        dina      => IL_L3PHIB_negPS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIB_negPS_2_B_V_readaddr,
        doutb     => IL_L3PHIB_negPS_2_B_V_dout,
        sync_nent => IL_L3PHIB_negPS_2_B_start,
        nent_o    => IL_L3PHIB_negPS_2_B_AV_dout_nent
      );

    IL_L3PHIB_negPS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIB_negPS_2_B_wea,
        addra     => IL_L3PHIB_negPS_2_B_writeaddr,
        dina      => IL_L3PHIB_negPS_2_B_din,
        wea_out       => IL_L3PHIB_negPS_2_B_wea_delay,
        addra_out     => IL_L3PHIB_negPS_2_B_writeaddr_delay,
        dina_out      => IL_L3PHIB_negPS_2_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHIB_negPS_2_B_start
      );

    IL_L3PHIC_negPS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHIC_negPS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHIC_negPS_2_B_wea_delay,
        addra     => IL_L3PHIC_negPS_2_B_writeaddr_delay,
        dina      => IL_L3PHIC_negPS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHIC_negPS_2_B_V_readaddr,
        doutb     => IL_L3PHIC_negPS_2_B_V_dout,
        sync_nent => IL_L3PHIC_negPS_2_B_start,
        nent_o    => IL_L3PHIC_negPS_2_B_AV_dout_nent
      );

    IL_L3PHIC_negPS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHIC_negPS_2_B_wea,
        addra     => IL_L3PHIC_negPS_2_B_writeaddr,
        dina      => IL_L3PHIC_negPS_2_B_din,
        wea_out       => IL_L3PHIC_negPS_2_B_wea_delay,
        addra_out     => IL_L3PHIC_negPS_2_B_writeaddr_delay,
        dina_out      => IL_L3PHIC_negPS_2_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHIC_negPS_2_B_start
      );

    IL_L3PHID_negPS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L3PHID_negPS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L3PHID_negPS_2_B_wea_delay,
        addra     => IL_L3PHID_negPS_2_B_writeaddr_delay,
        dina      => IL_L3PHID_negPS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L3PHID_negPS_2_B_V_readaddr,
        doutb     => IL_L3PHID_negPS_2_B_V_dout,
        sync_nent => IL_L3PHID_negPS_2_B_start,
        nent_o    => IL_L3PHID_negPS_2_B_AV_dout_nent
      );

    IL_L3PHID_negPS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L3PHID_negPS_2_B_wea,
        addra     => IL_L3PHID_negPS_2_B_writeaddr,
        dina      => IL_L3PHID_negPS_2_B_din,
        wea_out       => IL_L3PHID_negPS_2_B_wea_delay,
        addra_out     => IL_L3PHID_negPS_2_B_writeaddr_delay,
        dina_out      => IL_L3PHID_negPS_2_B_din_delay,
        done       => IR_done,
        start      => IL_L3PHID_negPS_2_B_start
      );

    IL_D4PHIA_negPS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIA_negPS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIA_negPS_2_A_wea_delay,
        addra     => IL_D4PHIA_negPS_2_A_writeaddr_delay,
        dina      => IL_D4PHIA_negPS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIA_negPS_2_A_V_readaddr,
        doutb     => IL_D4PHIA_negPS_2_A_V_dout,
        sync_nent => IL_D4PHIA_negPS_2_A_start,
        nent_o    => IL_D4PHIA_negPS_2_A_AV_dout_nent
      );

    IL_D4PHIA_negPS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIA_negPS_2_A_wea,
        addra     => IL_D4PHIA_negPS_2_A_writeaddr,
        dina      => IL_D4PHIA_negPS_2_A_din,
        wea_out       => IL_D4PHIA_negPS_2_A_wea_delay,
        addra_out     => IL_D4PHIA_negPS_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIA_negPS_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIA_negPS_2_A_start
      );

    IL_D4PHIB_negPS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_negPS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_negPS_2_A_wea_delay,
        addra     => IL_D4PHIB_negPS_2_A_writeaddr_delay,
        dina      => IL_D4PHIB_negPS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_negPS_2_A_V_readaddr,
        doutb     => IL_D4PHIB_negPS_2_A_V_dout,
        sync_nent => IL_D4PHIB_negPS_2_A_start,
        nent_o    => IL_D4PHIB_negPS_2_A_AV_dout_nent
      );

    IL_D4PHIB_negPS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_negPS_2_A_wea,
        addra     => IL_D4PHIB_negPS_2_A_writeaddr,
        dina      => IL_D4PHIB_negPS_2_A_din,
        wea_out       => IL_D4PHIB_negPS_2_A_wea_delay,
        addra_out     => IL_D4PHIB_negPS_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIB_negPS_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_negPS_2_A_start
      );

    IL_D4PHIB_negPS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_negPS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_negPS_2_B_wea_delay,
        addra     => IL_D4PHIB_negPS_2_B_writeaddr_delay,
        dina      => IL_D4PHIB_negPS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_negPS_2_B_V_readaddr,
        doutb     => IL_D4PHIB_negPS_2_B_V_dout,
        sync_nent => IL_D4PHIB_negPS_2_B_start,
        nent_o    => IL_D4PHIB_negPS_2_B_AV_dout_nent
      );

    IL_D4PHIB_negPS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_negPS_2_B_wea,
        addra     => IL_D4PHIB_negPS_2_B_writeaddr,
        dina      => IL_D4PHIB_negPS_2_B_din,
        wea_out       => IL_D4PHIB_negPS_2_B_wea_delay,
        addra_out     => IL_D4PHIB_negPS_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIB_negPS_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_negPS_2_B_start
      );

    IL_D4PHIC_negPS_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_negPS_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_negPS_2_A_wea_delay,
        addra     => IL_D4PHIC_negPS_2_A_writeaddr_delay,
        dina      => IL_D4PHIC_negPS_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_negPS_2_A_V_readaddr,
        doutb     => IL_D4PHIC_negPS_2_A_V_dout,
        sync_nent => IL_D4PHIC_negPS_2_A_start,
        nent_o    => IL_D4PHIC_negPS_2_A_AV_dout_nent
      );

    IL_D4PHIC_negPS_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_negPS_2_A_wea,
        addra     => IL_D4PHIC_negPS_2_A_writeaddr,
        dina      => IL_D4PHIC_negPS_2_A_din,
        wea_out       => IL_D4PHIC_negPS_2_A_wea_delay,
        addra_out     => IL_D4PHIC_negPS_2_A_writeaddr_delay,
        dina_out      => IL_D4PHIC_negPS_2_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_negPS_2_A_start
      );

    IL_D4PHIC_negPS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_negPS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_negPS_2_B_wea_delay,
        addra     => IL_D4PHIC_negPS_2_B_writeaddr_delay,
        dina      => IL_D4PHIC_negPS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_negPS_2_B_V_readaddr,
        doutb     => IL_D4PHIC_negPS_2_B_V_dout,
        sync_nent => IL_D4PHIC_negPS_2_B_start,
        nent_o    => IL_D4PHIC_negPS_2_B_AV_dout_nent
      );

    IL_D4PHIC_negPS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_negPS_2_B_wea,
        addra     => IL_D4PHIC_negPS_2_B_writeaddr,
        dina      => IL_D4PHIC_negPS_2_B_din,
        wea_out       => IL_D4PHIC_negPS_2_B_wea_delay,
        addra_out     => IL_D4PHIC_negPS_2_B_writeaddr_delay,
        dina_out      => IL_D4PHIC_negPS_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_negPS_2_B_start
      );

    IL_D4PHID_negPS_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHID_negPS_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHID_negPS_2_B_wea_delay,
        addra     => IL_D4PHID_negPS_2_B_writeaddr_delay,
        dina      => IL_D4PHID_negPS_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHID_negPS_2_B_V_readaddr,
        doutb     => IL_D4PHID_negPS_2_B_V_dout,
        sync_nent => IL_D4PHID_negPS_2_B_start,
        nent_o    => IL_D4PHID_negPS_2_B_AV_dout_nent
      );

    IL_D4PHID_negPS_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHID_negPS_2_B_wea,
        addra     => IL_D4PHID_negPS_2_B_writeaddr,
        dina      => IL_D4PHID_negPS_2_B_din,
        wea_out       => IL_D4PHID_negPS_2_B_wea_delay,
        addra_out     => IL_D4PHID_negPS_2_B_writeaddr_delay,
        dina_out      => IL_D4PHID_negPS_2_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHID_negPS_2_B_start
      );

    IL_L4PHIA_2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIA_2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIA_2S_1_A_wea_delay,
        addra     => IL_L4PHIA_2S_1_A_writeaddr_delay,
        dina      => IL_L4PHIA_2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIA_2S_1_A_V_readaddr,
        doutb     => IL_L4PHIA_2S_1_A_V_dout,
        sync_nent => IL_L4PHIA_2S_1_A_start,
        nent_o    => IL_L4PHIA_2S_1_A_AV_dout_nent
      );

    IL_L4PHIA_2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIA_2S_1_A_wea,
        addra     => IL_L4PHIA_2S_1_A_writeaddr,
        dina      => IL_L4PHIA_2S_1_A_din,
        wea_out       => IL_L4PHIA_2S_1_A_wea_delay,
        addra_out     => IL_L4PHIA_2S_1_A_writeaddr_delay,
        dina_out      => IL_L4PHIA_2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L4PHIA_2S_1_A_start
      );

    IL_L4PHIB_2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIB_2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIB_2S_1_A_wea_delay,
        addra     => IL_L4PHIB_2S_1_A_writeaddr_delay,
        dina      => IL_L4PHIB_2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIB_2S_1_A_V_readaddr,
        doutb     => IL_L4PHIB_2S_1_A_V_dout,
        sync_nent => IL_L4PHIB_2S_1_A_start,
        nent_o    => IL_L4PHIB_2S_1_A_AV_dout_nent
      );

    IL_L4PHIB_2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIB_2S_1_A_wea,
        addra     => IL_L4PHIB_2S_1_A_writeaddr,
        dina      => IL_L4PHIB_2S_1_A_din,
        wea_out       => IL_L4PHIB_2S_1_A_wea_delay,
        addra_out     => IL_L4PHIB_2S_1_A_writeaddr_delay,
        dina_out      => IL_L4PHIB_2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L4PHIB_2S_1_A_start
      );

    IL_L4PHIB_2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIB_2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIB_2S_1_B_wea_delay,
        addra     => IL_L4PHIB_2S_1_B_writeaddr_delay,
        dina      => IL_L4PHIB_2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIB_2S_1_B_V_readaddr,
        doutb     => IL_L4PHIB_2S_1_B_V_dout,
        sync_nent => IL_L4PHIB_2S_1_B_start,
        nent_o    => IL_L4PHIB_2S_1_B_AV_dout_nent
      );

    IL_L4PHIB_2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIB_2S_1_B_wea,
        addra     => IL_L4PHIB_2S_1_B_writeaddr,
        dina      => IL_L4PHIB_2S_1_B_din,
        wea_out       => IL_L4PHIB_2S_1_B_wea_delay,
        addra_out     => IL_L4PHIB_2S_1_B_writeaddr_delay,
        dina_out      => IL_L4PHIB_2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L4PHIB_2S_1_B_start
      );

    IL_L4PHIC_2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIC_2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIC_2S_1_A_wea_delay,
        addra     => IL_L4PHIC_2S_1_A_writeaddr_delay,
        dina      => IL_L4PHIC_2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIC_2S_1_A_V_readaddr,
        doutb     => IL_L4PHIC_2S_1_A_V_dout,
        sync_nent => IL_L4PHIC_2S_1_A_start,
        nent_o    => IL_L4PHIC_2S_1_A_AV_dout_nent
      );

    IL_L4PHIC_2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIC_2S_1_A_wea,
        addra     => IL_L4PHIC_2S_1_A_writeaddr,
        dina      => IL_L4PHIC_2S_1_A_din,
        wea_out       => IL_L4PHIC_2S_1_A_wea_delay,
        addra_out     => IL_L4PHIC_2S_1_A_writeaddr_delay,
        dina_out      => IL_L4PHIC_2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L4PHIC_2S_1_A_start
      );

    IL_L4PHIC_2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIC_2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIC_2S_1_B_wea_delay,
        addra     => IL_L4PHIC_2S_1_B_writeaddr_delay,
        dina      => IL_L4PHIC_2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIC_2S_1_B_V_readaddr,
        doutb     => IL_L4PHIC_2S_1_B_V_dout,
        sync_nent => IL_L4PHIC_2S_1_B_start,
        nent_o    => IL_L4PHIC_2S_1_B_AV_dout_nent
      );

    IL_L4PHIC_2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIC_2S_1_B_wea,
        addra     => IL_L4PHIC_2S_1_B_writeaddr,
        dina      => IL_L4PHIC_2S_1_B_din,
        wea_out       => IL_L4PHIC_2S_1_B_wea_delay,
        addra_out     => IL_L4PHIC_2S_1_B_writeaddr_delay,
        dina_out      => IL_L4PHIC_2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L4PHIC_2S_1_B_start
      );

    IL_L4PHID_2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHID_2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHID_2S_1_B_wea_delay,
        addra     => IL_L4PHID_2S_1_B_writeaddr_delay,
        dina      => IL_L4PHID_2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHID_2S_1_B_V_readaddr,
        doutb     => IL_L4PHID_2S_1_B_V_dout,
        sync_nent => IL_L4PHID_2S_1_B_start,
        nent_o    => IL_L4PHID_2S_1_B_AV_dout_nent
      );

    IL_L4PHID_2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHID_2S_1_B_wea,
        addra     => IL_L4PHID_2S_1_B_writeaddr,
        dina      => IL_L4PHID_2S_1_B_din,
        wea_out       => IL_L4PHID_2S_1_B_wea_delay,
        addra_out     => IL_L4PHID_2S_1_B_writeaddr_delay,
        dina_out      => IL_L4PHID_2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L4PHID_2S_1_B_start
      );

    IL_L5PHIA_2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIA_2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIA_2S_1_A_wea_delay,
        addra     => IL_L5PHIA_2S_1_A_writeaddr_delay,
        dina      => IL_L5PHIA_2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIA_2S_1_A_V_readaddr,
        doutb     => IL_L5PHIA_2S_1_A_V_dout,
        sync_nent => IL_L5PHIA_2S_1_A_start,
        nent_o    => IL_L5PHIA_2S_1_A_AV_dout_nent
      );

    IL_L5PHIA_2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIA_2S_1_A_wea,
        addra     => IL_L5PHIA_2S_1_A_writeaddr,
        dina      => IL_L5PHIA_2S_1_A_din,
        wea_out       => IL_L5PHIA_2S_1_A_wea_delay,
        addra_out     => IL_L5PHIA_2S_1_A_writeaddr_delay,
        dina_out      => IL_L5PHIA_2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIA_2S_1_A_start
      );

    IL_L5PHID_2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHID_2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHID_2S_1_B_wea_delay,
        addra     => IL_L5PHID_2S_1_B_writeaddr_delay,
        dina      => IL_L5PHID_2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHID_2S_1_B_V_readaddr,
        doutb     => IL_L5PHID_2S_1_B_V_dout,
        sync_nent => IL_L5PHID_2S_1_B_start,
        nent_o    => IL_L5PHID_2S_1_B_AV_dout_nent
      );

    IL_L5PHID_2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHID_2S_1_B_wea,
        addra     => IL_L5PHID_2S_1_B_writeaddr,
        dina      => IL_L5PHID_2S_1_B_din,
        wea_out       => IL_L5PHID_2S_1_B_wea_delay,
        addra_out     => IL_L5PHID_2S_1_B_writeaddr_delay,
        dina_out      => IL_L5PHID_2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHID_2S_1_B_start
      );

    IL_L5PHIA_2S_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIA_2S_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIA_2S_2_A_wea_delay,
        addra     => IL_L5PHIA_2S_2_A_writeaddr_delay,
        dina      => IL_L5PHIA_2S_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIA_2S_2_A_V_readaddr,
        doutb     => IL_L5PHIA_2S_2_A_V_dout,
        sync_nent => IL_L5PHIA_2S_2_A_start,
        nent_o    => IL_L5PHIA_2S_2_A_AV_dout_nent
      );

    IL_L5PHIA_2S_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIA_2S_2_A_wea,
        addra     => IL_L5PHIA_2S_2_A_writeaddr,
        dina      => IL_L5PHIA_2S_2_A_din,
        wea_out       => IL_L5PHIA_2S_2_A_wea_delay,
        addra_out     => IL_L5PHIA_2S_2_A_writeaddr_delay,
        dina_out      => IL_L5PHIA_2S_2_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIA_2S_2_A_start
      );

    IL_L5PHIB_2S_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIB_2S_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIB_2S_2_A_wea_delay,
        addra     => IL_L5PHIB_2S_2_A_writeaddr_delay,
        dina      => IL_L5PHIB_2S_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIB_2S_2_A_V_readaddr,
        doutb     => IL_L5PHIB_2S_2_A_V_dout,
        sync_nent => IL_L5PHIB_2S_2_A_start,
        nent_o    => IL_L5PHIB_2S_2_A_AV_dout_nent
      );

    IL_L5PHIB_2S_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIB_2S_2_A_wea,
        addra     => IL_L5PHIB_2S_2_A_writeaddr,
        dina      => IL_L5PHIB_2S_2_A_din,
        wea_out       => IL_L5PHIB_2S_2_A_wea_delay,
        addra_out     => IL_L5PHIB_2S_2_A_writeaddr_delay,
        dina_out      => IL_L5PHIB_2S_2_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIB_2S_2_A_start
      );

    IL_L5PHIB_2S_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIB_2S_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIB_2S_2_B_wea_delay,
        addra     => IL_L5PHIB_2S_2_B_writeaddr_delay,
        dina      => IL_L5PHIB_2S_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIB_2S_2_B_V_readaddr,
        doutb     => IL_L5PHIB_2S_2_B_V_dout,
        sync_nent => IL_L5PHIB_2S_2_B_start,
        nent_o    => IL_L5PHIB_2S_2_B_AV_dout_nent
      );

    IL_L5PHIB_2S_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIB_2S_2_B_wea,
        addra     => IL_L5PHIB_2S_2_B_writeaddr,
        dina      => IL_L5PHIB_2S_2_B_din,
        wea_out       => IL_L5PHIB_2S_2_B_wea_delay,
        addra_out     => IL_L5PHIB_2S_2_B_writeaddr_delay,
        dina_out      => IL_L5PHIB_2S_2_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHIB_2S_2_B_start
      );

    IL_L5PHIC_2S_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIC_2S_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIC_2S_2_A_wea_delay,
        addra     => IL_L5PHIC_2S_2_A_writeaddr_delay,
        dina      => IL_L5PHIC_2S_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIC_2S_2_A_V_readaddr,
        doutb     => IL_L5PHIC_2S_2_A_V_dout,
        sync_nent => IL_L5PHIC_2S_2_A_start,
        nent_o    => IL_L5PHIC_2S_2_A_AV_dout_nent
      );

    IL_L5PHIC_2S_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIC_2S_2_A_wea,
        addra     => IL_L5PHIC_2S_2_A_writeaddr,
        dina      => IL_L5PHIC_2S_2_A_din,
        wea_out       => IL_L5PHIC_2S_2_A_wea_delay,
        addra_out     => IL_L5PHIC_2S_2_A_writeaddr_delay,
        dina_out      => IL_L5PHIC_2S_2_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIC_2S_2_A_start
      );

    IL_L5PHIC_2S_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIC_2S_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIC_2S_2_B_wea_delay,
        addra     => IL_L5PHIC_2S_2_B_writeaddr_delay,
        dina      => IL_L5PHIC_2S_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIC_2S_2_B_V_readaddr,
        doutb     => IL_L5PHIC_2S_2_B_V_dout,
        sync_nent => IL_L5PHIC_2S_2_B_start,
        nent_o    => IL_L5PHIC_2S_2_B_AV_dout_nent
      );

    IL_L5PHIC_2S_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIC_2S_2_B_wea,
        addra     => IL_L5PHIC_2S_2_B_writeaddr,
        dina      => IL_L5PHIC_2S_2_B_din,
        wea_out       => IL_L5PHIC_2S_2_B_wea_delay,
        addra_out     => IL_L5PHIC_2S_2_B_writeaddr_delay,
        dina_out      => IL_L5PHIC_2S_2_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHIC_2S_2_B_start
      );

    IL_L5PHID_2S_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHID_2S_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHID_2S_2_B_wea_delay,
        addra     => IL_L5PHID_2S_2_B_writeaddr_delay,
        dina      => IL_L5PHID_2S_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHID_2S_2_B_V_readaddr,
        doutb     => IL_L5PHID_2S_2_B_V_dout,
        sync_nent => IL_L5PHID_2S_2_B_start,
        nent_o    => IL_L5PHID_2S_2_B_AV_dout_nent
      );

    IL_L5PHID_2S_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHID_2S_2_B_wea,
        addra     => IL_L5PHID_2S_2_B_writeaddr,
        dina      => IL_L5PHID_2S_2_B_din,
        wea_out       => IL_L5PHID_2S_2_B_wea_delay,
        addra_out     => IL_L5PHID_2S_2_B_writeaddr_delay,
        dina_out      => IL_L5PHID_2S_2_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHID_2S_2_B_start
      );

    IL_L6PHIA_2S_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIA_2S_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIA_2S_3_A_wea_delay,
        addra     => IL_L6PHIA_2S_3_A_writeaddr_delay,
        dina      => IL_L6PHIA_2S_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIA_2S_3_A_V_readaddr,
        doutb     => IL_L6PHIA_2S_3_A_V_dout,
        sync_nent => IL_L6PHIA_2S_3_A_start,
        nent_o    => IL_L6PHIA_2S_3_A_AV_dout_nent
      );

    IL_L6PHIA_2S_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIA_2S_3_A_wea,
        addra     => IL_L6PHIA_2S_3_A_writeaddr,
        dina      => IL_L6PHIA_2S_3_A_din,
        wea_out       => IL_L6PHIA_2S_3_A_wea_delay,
        addra_out     => IL_L6PHIA_2S_3_A_writeaddr_delay,
        dina_out      => IL_L6PHIA_2S_3_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIA_2S_3_A_start
      );

    IL_L6PHIB_2S_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIB_2S_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIB_2S_3_A_wea_delay,
        addra     => IL_L6PHIB_2S_3_A_writeaddr_delay,
        dina      => IL_L6PHIB_2S_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIB_2S_3_A_V_readaddr,
        doutb     => IL_L6PHIB_2S_3_A_V_dout,
        sync_nent => IL_L6PHIB_2S_3_A_start,
        nent_o    => IL_L6PHIB_2S_3_A_AV_dout_nent
      );

    IL_L6PHIB_2S_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIB_2S_3_A_wea,
        addra     => IL_L6PHIB_2S_3_A_writeaddr,
        dina      => IL_L6PHIB_2S_3_A_din,
        wea_out       => IL_L6PHIB_2S_3_A_wea_delay,
        addra_out     => IL_L6PHIB_2S_3_A_writeaddr_delay,
        dina_out      => IL_L6PHIB_2S_3_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIB_2S_3_A_start
      );

    IL_L6PHIC_2S_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIC_2S_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIC_2S_3_A_wea_delay,
        addra     => IL_L6PHIC_2S_3_A_writeaddr_delay,
        dina      => IL_L6PHIC_2S_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIC_2S_3_A_V_readaddr,
        doutb     => IL_L6PHIC_2S_3_A_V_dout,
        sync_nent => IL_L6PHIC_2S_3_A_start,
        nent_o    => IL_L6PHIC_2S_3_A_AV_dout_nent
      );

    IL_L6PHIC_2S_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIC_2S_3_A_wea,
        addra     => IL_L6PHIC_2S_3_A_writeaddr,
        dina      => IL_L6PHIC_2S_3_A_din,
        wea_out       => IL_L6PHIC_2S_3_A_wea_delay,
        addra_out     => IL_L6PHIC_2S_3_A_writeaddr_delay,
        dina_out      => IL_L6PHIC_2S_3_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIC_2S_3_A_start
      );

    IL_L6PHIC_2S_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIC_2S_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIC_2S_3_B_wea_delay,
        addra     => IL_L6PHIC_2S_3_B_writeaddr_delay,
        dina      => IL_L6PHIC_2S_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIC_2S_3_B_V_readaddr,
        doutb     => IL_L6PHIC_2S_3_B_V_dout,
        sync_nent => IL_L6PHIC_2S_3_B_start,
        nent_o    => IL_L6PHIC_2S_3_B_AV_dout_nent
      );

    IL_L6PHIC_2S_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIC_2S_3_B_wea,
        addra     => IL_L6PHIC_2S_3_B_writeaddr,
        dina      => IL_L6PHIC_2S_3_B_din,
        wea_out       => IL_L6PHIC_2S_3_B_wea_delay,
        addra_out     => IL_L6PHIC_2S_3_B_writeaddr_delay,
        dina_out      => IL_L6PHIC_2S_3_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHIC_2S_3_B_start
      );

    IL_L6PHID_2S_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHID_2S_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHID_2S_3_B_wea_delay,
        addra     => IL_L6PHID_2S_3_B_writeaddr_delay,
        dina      => IL_L6PHID_2S_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHID_2S_3_B_V_readaddr,
        doutb     => IL_L6PHID_2S_3_B_V_dout,
        sync_nent => IL_L6PHID_2S_3_B_start,
        nent_o    => IL_L6PHID_2S_3_B_AV_dout_nent
      );

    IL_L6PHID_2S_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHID_2S_3_B_wea,
        addra     => IL_L6PHID_2S_3_B_writeaddr,
        dina      => IL_L6PHID_2S_3_B_din,
        wea_out       => IL_L6PHID_2S_3_B_wea_delay,
        addra_out     => IL_L6PHID_2S_3_B_writeaddr_delay,
        dina_out      => IL_L6PHID_2S_3_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHID_2S_3_B_start
      );

    IL_L6PHIA_2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIA_2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIA_2S_4_A_wea_delay,
        addra     => IL_L6PHIA_2S_4_A_writeaddr_delay,
        dina      => IL_L6PHIA_2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIA_2S_4_A_V_readaddr,
        doutb     => IL_L6PHIA_2S_4_A_V_dout,
        sync_nent => IL_L6PHIA_2S_4_A_start,
        nent_o    => IL_L6PHIA_2S_4_A_AV_dout_nent
      );

    IL_L6PHIA_2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIA_2S_4_A_wea,
        addra     => IL_L6PHIA_2S_4_A_writeaddr,
        dina      => IL_L6PHIA_2S_4_A_din,
        wea_out       => IL_L6PHIA_2S_4_A_wea_delay,
        addra_out     => IL_L6PHIA_2S_4_A_writeaddr_delay,
        dina_out      => IL_L6PHIA_2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIA_2S_4_A_start
      );

    IL_L6PHIB_2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIB_2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIB_2S_4_A_wea_delay,
        addra     => IL_L6PHIB_2S_4_A_writeaddr_delay,
        dina      => IL_L6PHIB_2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIB_2S_4_A_V_readaddr,
        doutb     => IL_L6PHIB_2S_4_A_V_dout,
        sync_nent => IL_L6PHIB_2S_4_A_start,
        nent_o    => IL_L6PHIB_2S_4_A_AV_dout_nent
      );

    IL_L6PHIB_2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIB_2S_4_A_wea,
        addra     => IL_L6PHIB_2S_4_A_writeaddr,
        dina      => IL_L6PHIB_2S_4_A_din,
        wea_out       => IL_L6PHIB_2S_4_A_wea_delay,
        addra_out     => IL_L6PHIB_2S_4_A_writeaddr_delay,
        dina_out      => IL_L6PHIB_2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIB_2S_4_A_start
      );

    IL_L6PHIB_2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIB_2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIB_2S_4_B_wea_delay,
        addra     => IL_L6PHIB_2S_4_B_writeaddr_delay,
        dina      => IL_L6PHIB_2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIB_2S_4_B_V_readaddr,
        doutb     => IL_L6PHIB_2S_4_B_V_dout,
        sync_nent => IL_L6PHIB_2S_4_B_start,
        nent_o    => IL_L6PHIB_2S_4_B_AV_dout_nent
      );

    IL_L6PHIB_2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIB_2S_4_B_wea,
        addra     => IL_L6PHIB_2S_4_B_writeaddr,
        dina      => IL_L6PHIB_2S_4_B_din,
        wea_out       => IL_L6PHIB_2S_4_B_wea_delay,
        addra_out     => IL_L6PHIB_2S_4_B_writeaddr_delay,
        dina_out      => IL_L6PHIB_2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHIB_2S_4_B_start
      );

    IL_L6PHIC_2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIC_2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIC_2S_4_B_wea_delay,
        addra     => IL_L6PHIC_2S_4_B_writeaddr_delay,
        dina      => IL_L6PHIC_2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIC_2S_4_B_V_readaddr,
        doutb     => IL_L6PHIC_2S_4_B_V_dout,
        sync_nent => IL_L6PHIC_2S_4_B_start,
        nent_o    => IL_L6PHIC_2S_4_B_AV_dout_nent
      );

    IL_L6PHIC_2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIC_2S_4_B_wea,
        addra     => IL_L6PHIC_2S_4_B_writeaddr,
        dina      => IL_L6PHIC_2S_4_B_din,
        wea_out       => IL_L6PHIC_2S_4_B_wea_delay,
        addra_out     => IL_L6PHIC_2S_4_B_writeaddr_delay,
        dina_out      => IL_L6PHIC_2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHIC_2S_4_B_start
      );

    IL_L6PHID_2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHID_2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHID_2S_4_B_wea_delay,
        addra     => IL_L6PHID_2S_4_B_writeaddr_delay,
        dina      => IL_L6PHID_2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHID_2S_4_B_V_readaddr,
        doutb     => IL_L6PHID_2S_4_B_V_dout,
        sync_nent => IL_L6PHID_2S_4_B_start,
        nent_o    => IL_L6PHID_2S_4_B_AV_dout_nent
      );

    IL_L6PHID_2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHID_2S_4_B_wea,
        addra     => IL_L6PHID_2S_4_B_writeaddr,
        dina      => IL_L6PHID_2S_4_B_din,
        wea_out       => IL_L6PHID_2S_4_B_wea_delay,
        addra_out     => IL_L6PHID_2S_4_B_writeaddr_delay,
        dina_out      => IL_L6PHID_2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHID_2S_4_B_start
      );

    IL_D3PHIA_2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIA_2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIA_2S_4_A_wea_delay,
        addra     => IL_D3PHIA_2S_4_A_writeaddr_delay,
        dina      => IL_D3PHIA_2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIA_2S_4_A_V_readaddr,
        doutb     => IL_D3PHIA_2S_4_A_V_dout,
        sync_nent => IL_D3PHIA_2S_4_A_start,
        nent_o    => IL_D3PHIA_2S_4_A_AV_dout_nent
      );

    IL_D3PHIA_2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIA_2S_4_A_wea,
        addra     => IL_D3PHIA_2S_4_A_writeaddr,
        dina      => IL_D3PHIA_2S_4_A_din,
        wea_out       => IL_D3PHIA_2S_4_A_wea_delay,
        addra_out     => IL_D3PHIA_2S_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIA_2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIA_2S_4_A_start
      );

    IL_D3PHIB_2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_2S_4_A_wea_delay,
        addra     => IL_D3PHIB_2S_4_A_writeaddr_delay,
        dina      => IL_D3PHIB_2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_2S_4_A_V_readaddr,
        doutb     => IL_D3PHIB_2S_4_A_V_dout,
        sync_nent => IL_D3PHIB_2S_4_A_start,
        nent_o    => IL_D3PHIB_2S_4_A_AV_dout_nent
      );

    IL_D3PHIB_2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_2S_4_A_wea,
        addra     => IL_D3PHIB_2S_4_A_writeaddr,
        dina      => IL_D3PHIB_2S_4_A_din,
        wea_out       => IL_D3PHIB_2S_4_A_wea_delay,
        addra_out     => IL_D3PHIB_2S_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIB_2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_2S_4_A_start
      );

    IL_D3PHIB_2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_2S_4_B_wea_delay,
        addra     => IL_D3PHIB_2S_4_B_writeaddr_delay,
        dina      => IL_D3PHIB_2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_2S_4_B_V_readaddr,
        doutb     => IL_D3PHIB_2S_4_B_V_dout,
        sync_nent => IL_D3PHIB_2S_4_B_start,
        nent_o    => IL_D3PHIB_2S_4_B_AV_dout_nent
      );

    IL_D3PHIB_2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_2S_4_B_wea,
        addra     => IL_D3PHIB_2S_4_B_writeaddr,
        dina      => IL_D3PHIB_2S_4_B_din,
        wea_out       => IL_D3PHIB_2S_4_B_wea_delay,
        addra_out     => IL_D3PHIB_2S_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIB_2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_2S_4_B_start
      );

    IL_D3PHIC_2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_2S_4_A_wea_delay,
        addra     => IL_D3PHIC_2S_4_A_writeaddr_delay,
        dina      => IL_D3PHIC_2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_2S_4_A_V_readaddr,
        doutb     => IL_D3PHIC_2S_4_A_V_dout,
        sync_nent => IL_D3PHIC_2S_4_A_start,
        nent_o    => IL_D3PHIC_2S_4_A_AV_dout_nent
      );

    IL_D3PHIC_2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_2S_4_A_wea,
        addra     => IL_D3PHIC_2S_4_A_writeaddr,
        dina      => IL_D3PHIC_2S_4_A_din,
        wea_out       => IL_D3PHIC_2S_4_A_wea_delay,
        addra_out     => IL_D3PHIC_2S_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIC_2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_2S_4_A_start
      );

    IL_D3PHIC_2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_2S_4_B_wea_delay,
        addra     => IL_D3PHIC_2S_4_B_writeaddr_delay,
        dina      => IL_D3PHIC_2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_2S_4_B_V_readaddr,
        doutb     => IL_D3PHIC_2S_4_B_V_dout,
        sync_nent => IL_D3PHIC_2S_4_B_start,
        nent_o    => IL_D3PHIC_2S_4_B_AV_dout_nent
      );

    IL_D3PHIC_2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_2S_4_B_wea,
        addra     => IL_D3PHIC_2S_4_B_writeaddr,
        dina      => IL_D3PHIC_2S_4_B_din,
        wea_out       => IL_D3PHIC_2S_4_B_wea_delay,
        addra_out     => IL_D3PHIC_2S_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIC_2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_2S_4_B_start
      );

    IL_D3PHID_2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHID_2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHID_2S_4_B_wea_delay,
        addra     => IL_D3PHID_2S_4_B_writeaddr_delay,
        dina      => IL_D3PHID_2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHID_2S_4_B_V_readaddr,
        doutb     => IL_D3PHID_2S_4_B_V_dout,
        sync_nent => IL_D3PHID_2S_4_B_start,
        nent_o    => IL_D3PHID_2S_4_B_AV_dout_nent
      );

    IL_D3PHID_2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHID_2S_4_B_wea,
        addra     => IL_D3PHID_2S_4_B_writeaddr,
        dina      => IL_D3PHID_2S_4_B_din,
        wea_out       => IL_D3PHID_2S_4_B_wea_delay,
        addra_out     => IL_D3PHID_2S_4_B_writeaddr_delay,
        dina_out      => IL_D3PHID_2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHID_2S_4_B_start
      );

    IL_D1PHIA_2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIA_2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIA_2S_5_A_wea_delay,
        addra     => IL_D1PHIA_2S_5_A_writeaddr_delay,
        dina      => IL_D1PHIA_2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIA_2S_5_A_V_readaddr,
        doutb     => IL_D1PHIA_2S_5_A_V_dout,
        sync_nent => IL_D1PHIA_2S_5_A_start,
        nent_o    => IL_D1PHIA_2S_5_A_AV_dout_nent
      );

    IL_D1PHIA_2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIA_2S_5_A_wea,
        addra     => IL_D1PHIA_2S_5_A_writeaddr,
        dina      => IL_D1PHIA_2S_5_A_din,
        wea_out       => IL_D1PHIA_2S_5_A_wea_delay,
        addra_out     => IL_D1PHIA_2S_5_A_writeaddr_delay,
        dina_out      => IL_D1PHIA_2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIA_2S_5_A_start
      );

    IL_D1PHIB_2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_2S_5_A_wea_delay,
        addra     => IL_D1PHIB_2S_5_A_writeaddr_delay,
        dina      => IL_D1PHIB_2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_2S_5_A_V_readaddr,
        doutb     => IL_D1PHIB_2S_5_A_V_dout,
        sync_nent => IL_D1PHIB_2S_5_A_start,
        nent_o    => IL_D1PHIB_2S_5_A_AV_dout_nent
      );

    IL_D1PHIB_2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_2S_5_A_wea,
        addra     => IL_D1PHIB_2S_5_A_writeaddr,
        dina      => IL_D1PHIB_2S_5_A_din,
        wea_out       => IL_D1PHIB_2S_5_A_wea_delay,
        addra_out     => IL_D1PHIB_2S_5_A_writeaddr_delay,
        dina_out      => IL_D1PHIB_2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_2S_5_A_start
      );

    IL_D1PHIB_2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_2S_5_B_wea_delay,
        addra     => IL_D1PHIB_2S_5_B_writeaddr_delay,
        dina      => IL_D1PHIB_2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_2S_5_B_V_readaddr,
        doutb     => IL_D1PHIB_2S_5_B_V_dout,
        sync_nent => IL_D1PHIB_2S_5_B_start,
        nent_o    => IL_D1PHIB_2S_5_B_AV_dout_nent
      );

    IL_D1PHIB_2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_2S_5_B_wea,
        addra     => IL_D1PHIB_2S_5_B_writeaddr,
        dina      => IL_D1PHIB_2S_5_B_din,
        wea_out       => IL_D1PHIB_2S_5_B_wea_delay,
        addra_out     => IL_D1PHIB_2S_5_B_writeaddr_delay,
        dina_out      => IL_D1PHIB_2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_2S_5_B_start
      );

    IL_D1PHIC_2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_2S_5_A_wea_delay,
        addra     => IL_D1PHIC_2S_5_A_writeaddr_delay,
        dina      => IL_D1PHIC_2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_2S_5_A_V_readaddr,
        doutb     => IL_D1PHIC_2S_5_A_V_dout,
        sync_nent => IL_D1PHIC_2S_5_A_start,
        nent_o    => IL_D1PHIC_2S_5_A_AV_dout_nent
      );

    IL_D1PHIC_2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_2S_5_A_wea,
        addra     => IL_D1PHIC_2S_5_A_writeaddr,
        dina      => IL_D1PHIC_2S_5_A_din,
        wea_out       => IL_D1PHIC_2S_5_A_wea_delay,
        addra_out     => IL_D1PHIC_2S_5_A_writeaddr_delay,
        dina_out      => IL_D1PHIC_2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_2S_5_A_start
      );

    IL_D1PHIC_2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_2S_5_B_wea_delay,
        addra     => IL_D1PHIC_2S_5_B_writeaddr_delay,
        dina      => IL_D1PHIC_2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_2S_5_B_V_readaddr,
        doutb     => IL_D1PHIC_2S_5_B_V_dout,
        sync_nent => IL_D1PHIC_2S_5_B_start,
        nent_o    => IL_D1PHIC_2S_5_B_AV_dout_nent
      );

    IL_D1PHIC_2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_2S_5_B_wea,
        addra     => IL_D1PHIC_2S_5_B_writeaddr,
        dina      => IL_D1PHIC_2S_5_B_din,
        wea_out       => IL_D1PHIC_2S_5_B_wea_delay,
        addra_out     => IL_D1PHIC_2S_5_B_writeaddr_delay,
        dina_out      => IL_D1PHIC_2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_2S_5_B_start
      );

    IL_D1PHID_2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHID_2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHID_2S_5_B_wea_delay,
        addra     => IL_D1PHID_2S_5_B_writeaddr_delay,
        dina      => IL_D1PHID_2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHID_2S_5_B_V_readaddr,
        doutb     => IL_D1PHID_2S_5_B_V_dout,
        sync_nent => IL_D1PHID_2S_5_B_start,
        nent_o    => IL_D1PHID_2S_5_B_AV_dout_nent
      );

    IL_D1PHID_2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHID_2S_5_B_wea,
        addra     => IL_D1PHID_2S_5_B_writeaddr,
        dina      => IL_D1PHID_2S_5_B_din,
        wea_out       => IL_D1PHID_2S_5_B_wea_delay,
        addra_out     => IL_D1PHID_2S_5_B_writeaddr_delay,
        dina_out      => IL_D1PHID_2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHID_2S_5_B_start
      );

    IL_D4PHIA_2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIA_2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIA_2S_5_A_wea_delay,
        addra     => IL_D4PHIA_2S_5_A_writeaddr_delay,
        dina      => IL_D4PHIA_2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIA_2S_5_A_V_readaddr,
        doutb     => IL_D4PHIA_2S_5_A_V_dout,
        sync_nent => IL_D4PHIA_2S_5_A_start,
        nent_o    => IL_D4PHIA_2S_5_A_AV_dout_nent
      );

    IL_D4PHIA_2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIA_2S_5_A_wea,
        addra     => IL_D4PHIA_2S_5_A_writeaddr,
        dina      => IL_D4PHIA_2S_5_A_din,
        wea_out       => IL_D4PHIA_2S_5_A_wea_delay,
        addra_out     => IL_D4PHIA_2S_5_A_writeaddr_delay,
        dina_out      => IL_D4PHIA_2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIA_2S_5_A_start
      );

    IL_D4PHIB_2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_2S_5_A_wea_delay,
        addra     => IL_D4PHIB_2S_5_A_writeaddr_delay,
        dina      => IL_D4PHIB_2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_2S_5_A_V_readaddr,
        doutb     => IL_D4PHIB_2S_5_A_V_dout,
        sync_nent => IL_D4PHIB_2S_5_A_start,
        nent_o    => IL_D4PHIB_2S_5_A_AV_dout_nent
      );

    IL_D4PHIB_2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_2S_5_A_wea,
        addra     => IL_D4PHIB_2S_5_A_writeaddr,
        dina      => IL_D4PHIB_2S_5_A_din,
        wea_out       => IL_D4PHIB_2S_5_A_wea_delay,
        addra_out     => IL_D4PHIB_2S_5_A_writeaddr_delay,
        dina_out      => IL_D4PHIB_2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_2S_5_A_start
      );

    IL_D4PHIB_2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_2S_5_B_wea_delay,
        addra     => IL_D4PHIB_2S_5_B_writeaddr_delay,
        dina      => IL_D4PHIB_2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_2S_5_B_V_readaddr,
        doutb     => IL_D4PHIB_2S_5_B_V_dout,
        sync_nent => IL_D4PHIB_2S_5_B_start,
        nent_o    => IL_D4PHIB_2S_5_B_AV_dout_nent
      );

    IL_D4PHIB_2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_2S_5_B_wea,
        addra     => IL_D4PHIB_2S_5_B_writeaddr,
        dina      => IL_D4PHIB_2S_5_B_din,
        wea_out       => IL_D4PHIB_2S_5_B_wea_delay,
        addra_out     => IL_D4PHIB_2S_5_B_writeaddr_delay,
        dina_out      => IL_D4PHIB_2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_2S_5_B_start
      );

    IL_D4PHIC_2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_2S_5_A_wea_delay,
        addra     => IL_D4PHIC_2S_5_A_writeaddr_delay,
        dina      => IL_D4PHIC_2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_2S_5_A_V_readaddr,
        doutb     => IL_D4PHIC_2S_5_A_V_dout,
        sync_nent => IL_D4PHIC_2S_5_A_start,
        nent_o    => IL_D4PHIC_2S_5_A_AV_dout_nent
      );

    IL_D4PHIC_2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_2S_5_A_wea,
        addra     => IL_D4PHIC_2S_5_A_writeaddr,
        dina      => IL_D4PHIC_2S_5_A_din,
        wea_out       => IL_D4PHIC_2S_5_A_wea_delay,
        addra_out     => IL_D4PHIC_2S_5_A_writeaddr_delay,
        dina_out      => IL_D4PHIC_2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_2S_5_A_start
      );

    IL_D4PHIC_2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_2S_5_B_wea_delay,
        addra     => IL_D4PHIC_2S_5_B_writeaddr_delay,
        dina      => IL_D4PHIC_2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_2S_5_B_V_readaddr,
        doutb     => IL_D4PHIC_2S_5_B_V_dout,
        sync_nent => IL_D4PHIC_2S_5_B_start,
        nent_o    => IL_D4PHIC_2S_5_B_AV_dout_nent
      );

    IL_D4PHIC_2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_2S_5_B_wea,
        addra     => IL_D4PHIC_2S_5_B_writeaddr,
        dina      => IL_D4PHIC_2S_5_B_din,
        wea_out       => IL_D4PHIC_2S_5_B_wea_delay,
        addra_out     => IL_D4PHIC_2S_5_B_writeaddr_delay,
        dina_out      => IL_D4PHIC_2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_2S_5_B_start
      );

    IL_D4PHID_2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHID_2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHID_2S_5_B_wea_delay,
        addra     => IL_D4PHID_2S_5_B_writeaddr_delay,
        dina      => IL_D4PHID_2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHID_2S_5_B_V_readaddr,
        doutb     => IL_D4PHID_2S_5_B_V_dout,
        sync_nent => IL_D4PHID_2S_5_B_start,
        nent_o    => IL_D4PHID_2S_5_B_AV_dout_nent
      );

    IL_D4PHID_2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHID_2S_5_B_wea,
        addra     => IL_D4PHID_2S_5_B_writeaddr,
        dina      => IL_D4PHID_2S_5_B_din,
        wea_out       => IL_D4PHID_2S_5_B_wea_delay,
        addra_out     => IL_D4PHID_2S_5_B_writeaddr_delay,
        dina_out      => IL_D4PHID_2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHID_2S_5_B_start
      );

    IL_D2PHIA_2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_2S_6_A_wea_delay,
        addra     => IL_D2PHIA_2S_6_A_writeaddr_delay,
        dina      => IL_D2PHIA_2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_2S_6_A_V_readaddr,
        doutb     => IL_D2PHIA_2S_6_A_V_dout,
        sync_nent => IL_D2PHIA_2S_6_A_start,
        nent_o    => IL_D2PHIA_2S_6_A_AV_dout_nent
      );

    IL_D2PHIA_2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_2S_6_A_wea,
        addra     => IL_D2PHIA_2S_6_A_writeaddr,
        dina      => IL_D2PHIA_2S_6_A_din,
        wea_out       => IL_D2PHIA_2S_6_A_wea_delay,
        addra_out     => IL_D2PHIA_2S_6_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_2S_6_A_start
      );

    IL_D2PHIB_2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_2S_6_A_wea_delay,
        addra     => IL_D2PHIB_2S_6_A_writeaddr_delay,
        dina      => IL_D2PHIB_2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_2S_6_A_V_readaddr,
        doutb     => IL_D2PHIB_2S_6_A_V_dout,
        sync_nent => IL_D2PHIB_2S_6_A_start,
        nent_o    => IL_D2PHIB_2S_6_A_AV_dout_nent
      );

    IL_D2PHIB_2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_2S_6_A_wea,
        addra     => IL_D2PHIB_2S_6_A_writeaddr,
        dina      => IL_D2PHIB_2S_6_A_din,
        wea_out       => IL_D2PHIB_2S_6_A_wea_delay,
        addra_out     => IL_D2PHIB_2S_6_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_2S_6_A_start
      );

    IL_D2PHIB_2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_2S_6_B_wea_delay,
        addra     => IL_D2PHIB_2S_6_B_writeaddr_delay,
        dina      => IL_D2PHIB_2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_2S_6_B_V_readaddr,
        doutb     => IL_D2PHIB_2S_6_B_V_dout,
        sync_nent => IL_D2PHIB_2S_6_B_start,
        nent_o    => IL_D2PHIB_2S_6_B_AV_dout_nent
      );

    IL_D2PHIB_2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_2S_6_B_wea,
        addra     => IL_D2PHIB_2S_6_B_writeaddr,
        dina      => IL_D2PHIB_2S_6_B_din,
        wea_out       => IL_D2PHIB_2S_6_B_wea_delay,
        addra_out     => IL_D2PHIB_2S_6_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_2S_6_B_start
      );

    IL_D2PHIC_2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_2S_6_A_wea_delay,
        addra     => IL_D2PHIC_2S_6_A_writeaddr_delay,
        dina      => IL_D2PHIC_2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_2S_6_A_V_readaddr,
        doutb     => IL_D2PHIC_2S_6_A_V_dout,
        sync_nent => IL_D2PHIC_2S_6_A_start,
        nent_o    => IL_D2PHIC_2S_6_A_AV_dout_nent
      );

    IL_D2PHIC_2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_2S_6_A_wea,
        addra     => IL_D2PHIC_2S_6_A_writeaddr,
        dina      => IL_D2PHIC_2S_6_A_din,
        wea_out       => IL_D2PHIC_2S_6_A_wea_delay,
        addra_out     => IL_D2PHIC_2S_6_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_2S_6_A_start
      );

    IL_D2PHIC_2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_2S_6_B_wea_delay,
        addra     => IL_D2PHIC_2S_6_B_writeaddr_delay,
        dina      => IL_D2PHIC_2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_2S_6_B_V_readaddr,
        doutb     => IL_D2PHIC_2S_6_B_V_dout,
        sync_nent => IL_D2PHIC_2S_6_B_start,
        nent_o    => IL_D2PHIC_2S_6_B_AV_dout_nent
      );

    IL_D2PHIC_2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_2S_6_B_wea,
        addra     => IL_D2PHIC_2S_6_B_writeaddr,
        dina      => IL_D2PHIC_2S_6_B_din,
        wea_out       => IL_D2PHIC_2S_6_B_wea_delay,
        addra_out     => IL_D2PHIC_2S_6_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_2S_6_B_start
      );

    IL_D2PHID_2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_2S_6_B_wea_delay,
        addra     => IL_D2PHID_2S_6_B_writeaddr_delay,
        dina      => IL_D2PHID_2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_2S_6_B_V_readaddr,
        doutb     => IL_D2PHID_2S_6_B_V_dout,
        sync_nent => IL_D2PHID_2S_6_B_start,
        nent_o    => IL_D2PHID_2S_6_B_AV_dout_nent
      );

    IL_D2PHID_2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_2S_6_B_wea,
        addra     => IL_D2PHID_2S_6_B_writeaddr,
        dina      => IL_D2PHID_2S_6_B_din,
        wea_out       => IL_D2PHID_2S_6_B_wea_delay,
        addra_out     => IL_D2PHID_2S_6_B_writeaddr_delay,
        dina_out      => IL_D2PHID_2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_2S_6_B_start
      );

    IL_D5PHIA_2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIA_2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIA_2S_6_A_wea_delay,
        addra     => IL_D5PHIA_2S_6_A_writeaddr_delay,
        dina      => IL_D5PHIA_2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIA_2S_6_A_V_readaddr,
        doutb     => IL_D5PHIA_2S_6_A_V_dout,
        sync_nent => IL_D5PHIA_2S_6_A_start,
        nent_o    => IL_D5PHIA_2S_6_A_AV_dout_nent
      );

    IL_D5PHIA_2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIA_2S_6_A_wea,
        addra     => IL_D5PHIA_2S_6_A_writeaddr,
        dina      => IL_D5PHIA_2S_6_A_din,
        wea_out       => IL_D5PHIA_2S_6_A_wea_delay,
        addra_out     => IL_D5PHIA_2S_6_A_writeaddr_delay,
        dina_out      => IL_D5PHIA_2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIA_2S_6_A_start
      );

    IL_D5PHIB_2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_2S_6_A_wea_delay,
        addra     => IL_D5PHIB_2S_6_A_writeaddr_delay,
        dina      => IL_D5PHIB_2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_2S_6_A_V_readaddr,
        doutb     => IL_D5PHIB_2S_6_A_V_dout,
        sync_nent => IL_D5PHIB_2S_6_A_start,
        nent_o    => IL_D5PHIB_2S_6_A_AV_dout_nent
      );

    IL_D5PHIB_2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_2S_6_A_wea,
        addra     => IL_D5PHIB_2S_6_A_writeaddr,
        dina      => IL_D5PHIB_2S_6_A_din,
        wea_out       => IL_D5PHIB_2S_6_A_wea_delay,
        addra_out     => IL_D5PHIB_2S_6_A_writeaddr_delay,
        dina_out      => IL_D5PHIB_2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_2S_6_A_start
      );

    IL_D5PHIB_2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_2S_6_B_wea_delay,
        addra     => IL_D5PHIB_2S_6_B_writeaddr_delay,
        dina      => IL_D5PHIB_2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_2S_6_B_V_readaddr,
        doutb     => IL_D5PHIB_2S_6_B_V_dout,
        sync_nent => IL_D5PHIB_2S_6_B_start,
        nent_o    => IL_D5PHIB_2S_6_B_AV_dout_nent
      );

    IL_D5PHIB_2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_2S_6_B_wea,
        addra     => IL_D5PHIB_2S_6_B_writeaddr,
        dina      => IL_D5PHIB_2S_6_B_din,
        wea_out       => IL_D5PHIB_2S_6_B_wea_delay,
        addra_out     => IL_D5PHIB_2S_6_B_writeaddr_delay,
        dina_out      => IL_D5PHIB_2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_2S_6_B_start
      );

    IL_D5PHIC_2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_2S_6_A_wea_delay,
        addra     => IL_D5PHIC_2S_6_A_writeaddr_delay,
        dina      => IL_D5PHIC_2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_2S_6_A_V_readaddr,
        doutb     => IL_D5PHIC_2S_6_A_V_dout,
        sync_nent => IL_D5PHIC_2S_6_A_start,
        nent_o    => IL_D5PHIC_2S_6_A_AV_dout_nent
      );

    IL_D5PHIC_2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_2S_6_A_wea,
        addra     => IL_D5PHIC_2S_6_A_writeaddr,
        dina      => IL_D5PHIC_2S_6_A_din,
        wea_out       => IL_D5PHIC_2S_6_A_wea_delay,
        addra_out     => IL_D5PHIC_2S_6_A_writeaddr_delay,
        dina_out      => IL_D5PHIC_2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_2S_6_A_start
      );

    IL_D5PHIC_2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_2S_6_B_wea_delay,
        addra     => IL_D5PHIC_2S_6_B_writeaddr_delay,
        dina      => IL_D5PHIC_2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_2S_6_B_V_readaddr,
        doutb     => IL_D5PHIC_2S_6_B_V_dout,
        sync_nent => IL_D5PHIC_2S_6_B_start,
        nent_o    => IL_D5PHIC_2S_6_B_AV_dout_nent
      );

    IL_D5PHIC_2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_2S_6_B_wea,
        addra     => IL_D5PHIC_2S_6_B_writeaddr,
        dina      => IL_D5PHIC_2S_6_B_din,
        wea_out       => IL_D5PHIC_2S_6_B_wea_delay,
        addra_out     => IL_D5PHIC_2S_6_B_writeaddr_delay,
        dina_out      => IL_D5PHIC_2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_2S_6_B_start
      );

    IL_D5PHID_2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHID_2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHID_2S_6_B_wea_delay,
        addra     => IL_D5PHID_2S_6_B_writeaddr_delay,
        dina      => IL_D5PHID_2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHID_2S_6_B_V_readaddr,
        doutb     => IL_D5PHID_2S_6_B_V_dout,
        sync_nent => IL_D5PHID_2S_6_B_start,
        nent_o    => IL_D5PHID_2S_6_B_AV_dout_nent
      );

    IL_D5PHID_2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHID_2S_6_B_wea,
        addra     => IL_D5PHID_2S_6_B_writeaddr,
        dina      => IL_D5PHID_2S_6_B_din,
        wea_out       => IL_D5PHID_2S_6_B_wea_delay,
        addra_out     => IL_D5PHID_2S_6_B_writeaddr_delay,
        dina_out      => IL_D5PHID_2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHID_2S_6_B_start
      );

    IL_L4PHIA_neg2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIA_neg2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIA_neg2S_1_A_wea_delay,
        addra     => IL_L4PHIA_neg2S_1_A_writeaddr_delay,
        dina      => IL_L4PHIA_neg2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIA_neg2S_1_A_V_readaddr,
        doutb     => IL_L4PHIA_neg2S_1_A_V_dout,
        sync_nent => IL_L4PHIA_neg2S_1_A_start,
        nent_o    => IL_L4PHIA_neg2S_1_A_AV_dout_nent
      );

    IL_L4PHIA_neg2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIA_neg2S_1_A_wea,
        addra     => IL_L4PHIA_neg2S_1_A_writeaddr,
        dina      => IL_L4PHIA_neg2S_1_A_din,
        wea_out       => IL_L4PHIA_neg2S_1_A_wea_delay,
        addra_out     => IL_L4PHIA_neg2S_1_A_writeaddr_delay,
        dina_out      => IL_L4PHIA_neg2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L4PHIA_neg2S_1_A_start
      );

    IL_L4PHIB_neg2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIB_neg2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIB_neg2S_1_A_wea_delay,
        addra     => IL_L4PHIB_neg2S_1_A_writeaddr_delay,
        dina      => IL_L4PHIB_neg2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIB_neg2S_1_A_V_readaddr,
        doutb     => IL_L4PHIB_neg2S_1_A_V_dout,
        sync_nent => IL_L4PHIB_neg2S_1_A_start,
        nent_o    => IL_L4PHIB_neg2S_1_A_AV_dout_nent
      );

    IL_L4PHIB_neg2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIB_neg2S_1_A_wea,
        addra     => IL_L4PHIB_neg2S_1_A_writeaddr,
        dina      => IL_L4PHIB_neg2S_1_A_din,
        wea_out       => IL_L4PHIB_neg2S_1_A_wea_delay,
        addra_out     => IL_L4PHIB_neg2S_1_A_writeaddr_delay,
        dina_out      => IL_L4PHIB_neg2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L4PHIB_neg2S_1_A_start
      );

    IL_L4PHIB_neg2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIB_neg2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIB_neg2S_1_B_wea_delay,
        addra     => IL_L4PHIB_neg2S_1_B_writeaddr_delay,
        dina      => IL_L4PHIB_neg2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIB_neg2S_1_B_V_readaddr,
        doutb     => IL_L4PHIB_neg2S_1_B_V_dout,
        sync_nent => IL_L4PHIB_neg2S_1_B_start,
        nent_o    => IL_L4PHIB_neg2S_1_B_AV_dout_nent
      );

    IL_L4PHIB_neg2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIB_neg2S_1_B_wea,
        addra     => IL_L4PHIB_neg2S_1_B_writeaddr,
        dina      => IL_L4PHIB_neg2S_1_B_din,
        wea_out       => IL_L4PHIB_neg2S_1_B_wea_delay,
        addra_out     => IL_L4PHIB_neg2S_1_B_writeaddr_delay,
        dina_out      => IL_L4PHIB_neg2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L4PHIB_neg2S_1_B_start
      );

    IL_L4PHIC_neg2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIC_neg2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIC_neg2S_1_A_wea_delay,
        addra     => IL_L4PHIC_neg2S_1_A_writeaddr_delay,
        dina      => IL_L4PHIC_neg2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIC_neg2S_1_A_V_readaddr,
        doutb     => IL_L4PHIC_neg2S_1_A_V_dout,
        sync_nent => IL_L4PHIC_neg2S_1_A_start,
        nent_o    => IL_L4PHIC_neg2S_1_A_AV_dout_nent
      );

    IL_L4PHIC_neg2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIC_neg2S_1_A_wea,
        addra     => IL_L4PHIC_neg2S_1_A_writeaddr,
        dina      => IL_L4PHIC_neg2S_1_A_din,
        wea_out       => IL_L4PHIC_neg2S_1_A_wea_delay,
        addra_out     => IL_L4PHIC_neg2S_1_A_writeaddr_delay,
        dina_out      => IL_L4PHIC_neg2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L4PHIC_neg2S_1_A_start
      );

    IL_L4PHIC_neg2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHIC_neg2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHIC_neg2S_1_B_wea_delay,
        addra     => IL_L4PHIC_neg2S_1_B_writeaddr_delay,
        dina      => IL_L4PHIC_neg2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHIC_neg2S_1_B_V_readaddr,
        doutb     => IL_L4PHIC_neg2S_1_B_V_dout,
        sync_nent => IL_L4PHIC_neg2S_1_B_start,
        nent_o    => IL_L4PHIC_neg2S_1_B_AV_dout_nent
      );

    IL_L4PHIC_neg2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHIC_neg2S_1_B_wea,
        addra     => IL_L4PHIC_neg2S_1_B_writeaddr,
        dina      => IL_L4PHIC_neg2S_1_B_din,
        wea_out       => IL_L4PHIC_neg2S_1_B_wea_delay,
        addra_out     => IL_L4PHIC_neg2S_1_B_writeaddr_delay,
        dina_out      => IL_L4PHIC_neg2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L4PHIC_neg2S_1_B_start
      );

    IL_L4PHID_neg2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L4PHID_neg2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L4PHID_neg2S_1_B_wea_delay,
        addra     => IL_L4PHID_neg2S_1_B_writeaddr_delay,
        dina      => IL_L4PHID_neg2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L4PHID_neg2S_1_B_V_readaddr,
        doutb     => IL_L4PHID_neg2S_1_B_V_dout,
        sync_nent => IL_L4PHID_neg2S_1_B_start,
        nent_o    => IL_L4PHID_neg2S_1_B_AV_dout_nent
      );

    IL_L4PHID_neg2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L4PHID_neg2S_1_B_wea,
        addra     => IL_L4PHID_neg2S_1_B_writeaddr,
        dina      => IL_L4PHID_neg2S_1_B_din,
        wea_out       => IL_L4PHID_neg2S_1_B_wea_delay,
        addra_out     => IL_L4PHID_neg2S_1_B_writeaddr_delay,
        dina_out      => IL_L4PHID_neg2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L4PHID_neg2S_1_B_start
      );

    IL_L5PHIA_neg2S_1_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIA_neg2S_1_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIA_neg2S_1_A_wea_delay,
        addra     => IL_L5PHIA_neg2S_1_A_writeaddr_delay,
        dina      => IL_L5PHIA_neg2S_1_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIA_neg2S_1_A_V_readaddr,
        doutb     => IL_L5PHIA_neg2S_1_A_V_dout,
        sync_nent => IL_L5PHIA_neg2S_1_A_start,
        nent_o    => IL_L5PHIA_neg2S_1_A_AV_dout_nent
      );

    IL_L5PHIA_neg2S_1_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIA_neg2S_1_A_wea,
        addra     => IL_L5PHIA_neg2S_1_A_writeaddr,
        dina      => IL_L5PHIA_neg2S_1_A_din,
        wea_out       => IL_L5PHIA_neg2S_1_A_wea_delay,
        addra_out     => IL_L5PHIA_neg2S_1_A_writeaddr_delay,
        dina_out      => IL_L5PHIA_neg2S_1_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIA_neg2S_1_A_start
      );

    IL_L5PHID_neg2S_1_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHID_neg2S_1_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHID_neg2S_1_B_wea_delay,
        addra     => IL_L5PHID_neg2S_1_B_writeaddr_delay,
        dina      => IL_L5PHID_neg2S_1_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHID_neg2S_1_B_V_readaddr,
        doutb     => IL_L5PHID_neg2S_1_B_V_dout,
        sync_nent => IL_L5PHID_neg2S_1_B_start,
        nent_o    => IL_L5PHID_neg2S_1_B_AV_dout_nent
      );

    IL_L5PHID_neg2S_1_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHID_neg2S_1_B_wea,
        addra     => IL_L5PHID_neg2S_1_B_writeaddr,
        dina      => IL_L5PHID_neg2S_1_B_din,
        wea_out       => IL_L5PHID_neg2S_1_B_wea_delay,
        addra_out     => IL_L5PHID_neg2S_1_B_writeaddr_delay,
        dina_out      => IL_L5PHID_neg2S_1_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHID_neg2S_1_B_start
      );

    IL_L5PHIA_neg2S_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIA_neg2S_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIA_neg2S_2_A_wea_delay,
        addra     => IL_L5PHIA_neg2S_2_A_writeaddr_delay,
        dina      => IL_L5PHIA_neg2S_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIA_neg2S_2_A_V_readaddr,
        doutb     => IL_L5PHIA_neg2S_2_A_V_dout,
        sync_nent => IL_L5PHIA_neg2S_2_A_start,
        nent_o    => IL_L5PHIA_neg2S_2_A_AV_dout_nent
      );

    IL_L5PHIA_neg2S_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIA_neg2S_2_A_wea,
        addra     => IL_L5PHIA_neg2S_2_A_writeaddr,
        dina      => IL_L5PHIA_neg2S_2_A_din,
        wea_out       => IL_L5PHIA_neg2S_2_A_wea_delay,
        addra_out     => IL_L5PHIA_neg2S_2_A_writeaddr_delay,
        dina_out      => IL_L5PHIA_neg2S_2_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIA_neg2S_2_A_start
      );

    IL_L5PHIB_neg2S_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIB_neg2S_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIB_neg2S_2_A_wea_delay,
        addra     => IL_L5PHIB_neg2S_2_A_writeaddr_delay,
        dina      => IL_L5PHIB_neg2S_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIB_neg2S_2_A_V_readaddr,
        doutb     => IL_L5PHIB_neg2S_2_A_V_dout,
        sync_nent => IL_L5PHIB_neg2S_2_A_start,
        nent_o    => IL_L5PHIB_neg2S_2_A_AV_dout_nent
      );

    IL_L5PHIB_neg2S_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIB_neg2S_2_A_wea,
        addra     => IL_L5PHIB_neg2S_2_A_writeaddr,
        dina      => IL_L5PHIB_neg2S_2_A_din,
        wea_out       => IL_L5PHIB_neg2S_2_A_wea_delay,
        addra_out     => IL_L5PHIB_neg2S_2_A_writeaddr_delay,
        dina_out      => IL_L5PHIB_neg2S_2_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIB_neg2S_2_A_start
      );

    IL_L5PHIB_neg2S_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIB_neg2S_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIB_neg2S_2_B_wea_delay,
        addra     => IL_L5PHIB_neg2S_2_B_writeaddr_delay,
        dina      => IL_L5PHIB_neg2S_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIB_neg2S_2_B_V_readaddr,
        doutb     => IL_L5PHIB_neg2S_2_B_V_dout,
        sync_nent => IL_L5PHIB_neg2S_2_B_start,
        nent_o    => IL_L5PHIB_neg2S_2_B_AV_dout_nent
      );

    IL_L5PHIB_neg2S_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIB_neg2S_2_B_wea,
        addra     => IL_L5PHIB_neg2S_2_B_writeaddr,
        dina      => IL_L5PHIB_neg2S_2_B_din,
        wea_out       => IL_L5PHIB_neg2S_2_B_wea_delay,
        addra_out     => IL_L5PHIB_neg2S_2_B_writeaddr_delay,
        dina_out      => IL_L5PHIB_neg2S_2_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHIB_neg2S_2_B_start
      );

    IL_L5PHIC_neg2S_2_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIC_neg2S_2_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIC_neg2S_2_A_wea_delay,
        addra     => IL_L5PHIC_neg2S_2_A_writeaddr_delay,
        dina      => IL_L5PHIC_neg2S_2_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIC_neg2S_2_A_V_readaddr,
        doutb     => IL_L5PHIC_neg2S_2_A_V_dout,
        sync_nent => IL_L5PHIC_neg2S_2_A_start,
        nent_o    => IL_L5PHIC_neg2S_2_A_AV_dout_nent
      );

    IL_L5PHIC_neg2S_2_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIC_neg2S_2_A_wea,
        addra     => IL_L5PHIC_neg2S_2_A_writeaddr,
        dina      => IL_L5PHIC_neg2S_2_A_din,
        wea_out       => IL_L5PHIC_neg2S_2_A_wea_delay,
        addra_out     => IL_L5PHIC_neg2S_2_A_writeaddr_delay,
        dina_out      => IL_L5PHIC_neg2S_2_A_din_delay,
        done       => IR_done,
        start      => IL_L5PHIC_neg2S_2_A_start
      );

    IL_L5PHIC_neg2S_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHIC_neg2S_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHIC_neg2S_2_B_wea_delay,
        addra     => IL_L5PHIC_neg2S_2_B_writeaddr_delay,
        dina      => IL_L5PHIC_neg2S_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHIC_neg2S_2_B_V_readaddr,
        doutb     => IL_L5PHIC_neg2S_2_B_V_dout,
        sync_nent => IL_L5PHIC_neg2S_2_B_start,
        nent_o    => IL_L5PHIC_neg2S_2_B_AV_dout_nent
      );

    IL_L5PHIC_neg2S_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHIC_neg2S_2_B_wea,
        addra     => IL_L5PHIC_neg2S_2_B_writeaddr,
        dina      => IL_L5PHIC_neg2S_2_B_din,
        wea_out       => IL_L5PHIC_neg2S_2_B_wea_delay,
        addra_out     => IL_L5PHIC_neg2S_2_B_writeaddr_delay,
        dina_out      => IL_L5PHIC_neg2S_2_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHIC_neg2S_2_B_start
      );

    IL_L5PHID_neg2S_2_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L5PHID_neg2S_2_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L5PHID_neg2S_2_B_wea_delay,
        addra     => IL_L5PHID_neg2S_2_B_writeaddr_delay,
        dina      => IL_L5PHID_neg2S_2_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L5PHID_neg2S_2_B_V_readaddr,
        doutb     => IL_L5PHID_neg2S_2_B_V_dout,
        sync_nent => IL_L5PHID_neg2S_2_B_start,
        nent_o    => IL_L5PHID_neg2S_2_B_AV_dout_nent
      );

    IL_L5PHID_neg2S_2_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L5PHID_neg2S_2_B_wea,
        addra     => IL_L5PHID_neg2S_2_B_writeaddr,
        dina      => IL_L5PHID_neg2S_2_B_din,
        wea_out       => IL_L5PHID_neg2S_2_B_wea_delay,
        addra_out     => IL_L5PHID_neg2S_2_B_writeaddr_delay,
        dina_out      => IL_L5PHID_neg2S_2_B_din_delay,
        done       => IR_done,
        start      => IL_L5PHID_neg2S_2_B_start
      );

    IL_L6PHIA_neg2S_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIA_neg2S_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIA_neg2S_3_A_wea_delay,
        addra     => IL_L6PHIA_neg2S_3_A_writeaddr_delay,
        dina      => IL_L6PHIA_neg2S_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIA_neg2S_3_A_V_readaddr,
        doutb     => IL_L6PHIA_neg2S_3_A_V_dout,
        sync_nent => IL_L6PHIA_neg2S_3_A_start,
        nent_o    => IL_L6PHIA_neg2S_3_A_AV_dout_nent
      );

    IL_L6PHIA_neg2S_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIA_neg2S_3_A_wea,
        addra     => IL_L6PHIA_neg2S_3_A_writeaddr,
        dina      => IL_L6PHIA_neg2S_3_A_din,
        wea_out       => IL_L6PHIA_neg2S_3_A_wea_delay,
        addra_out     => IL_L6PHIA_neg2S_3_A_writeaddr_delay,
        dina_out      => IL_L6PHIA_neg2S_3_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIA_neg2S_3_A_start
      );

    IL_L6PHIB_neg2S_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIB_neg2S_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIB_neg2S_3_A_wea_delay,
        addra     => IL_L6PHIB_neg2S_3_A_writeaddr_delay,
        dina      => IL_L6PHIB_neg2S_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIB_neg2S_3_A_V_readaddr,
        doutb     => IL_L6PHIB_neg2S_3_A_V_dout,
        sync_nent => IL_L6PHIB_neg2S_3_A_start,
        nent_o    => IL_L6PHIB_neg2S_3_A_AV_dout_nent
      );

    IL_L6PHIB_neg2S_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIB_neg2S_3_A_wea,
        addra     => IL_L6PHIB_neg2S_3_A_writeaddr,
        dina      => IL_L6PHIB_neg2S_3_A_din,
        wea_out       => IL_L6PHIB_neg2S_3_A_wea_delay,
        addra_out     => IL_L6PHIB_neg2S_3_A_writeaddr_delay,
        dina_out      => IL_L6PHIB_neg2S_3_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIB_neg2S_3_A_start
      );

    IL_L6PHIC_neg2S_3_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIC_neg2S_3_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIC_neg2S_3_A_wea_delay,
        addra     => IL_L6PHIC_neg2S_3_A_writeaddr_delay,
        dina      => IL_L6PHIC_neg2S_3_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIC_neg2S_3_A_V_readaddr,
        doutb     => IL_L6PHIC_neg2S_3_A_V_dout,
        sync_nent => IL_L6PHIC_neg2S_3_A_start,
        nent_o    => IL_L6PHIC_neg2S_3_A_AV_dout_nent
      );

    IL_L6PHIC_neg2S_3_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIC_neg2S_3_A_wea,
        addra     => IL_L6PHIC_neg2S_3_A_writeaddr,
        dina      => IL_L6PHIC_neg2S_3_A_din,
        wea_out       => IL_L6PHIC_neg2S_3_A_wea_delay,
        addra_out     => IL_L6PHIC_neg2S_3_A_writeaddr_delay,
        dina_out      => IL_L6PHIC_neg2S_3_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIC_neg2S_3_A_start
      );

    IL_L6PHIC_neg2S_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIC_neg2S_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIC_neg2S_3_B_wea_delay,
        addra     => IL_L6PHIC_neg2S_3_B_writeaddr_delay,
        dina      => IL_L6PHIC_neg2S_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIC_neg2S_3_B_V_readaddr,
        doutb     => IL_L6PHIC_neg2S_3_B_V_dout,
        sync_nent => IL_L6PHIC_neg2S_3_B_start,
        nent_o    => IL_L6PHIC_neg2S_3_B_AV_dout_nent
      );

    IL_L6PHIC_neg2S_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIC_neg2S_3_B_wea,
        addra     => IL_L6PHIC_neg2S_3_B_writeaddr,
        dina      => IL_L6PHIC_neg2S_3_B_din,
        wea_out       => IL_L6PHIC_neg2S_3_B_wea_delay,
        addra_out     => IL_L6PHIC_neg2S_3_B_writeaddr_delay,
        dina_out      => IL_L6PHIC_neg2S_3_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHIC_neg2S_3_B_start
      );

    IL_L6PHID_neg2S_3_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHID_neg2S_3_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHID_neg2S_3_B_wea_delay,
        addra     => IL_L6PHID_neg2S_3_B_writeaddr_delay,
        dina      => IL_L6PHID_neg2S_3_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHID_neg2S_3_B_V_readaddr,
        doutb     => IL_L6PHID_neg2S_3_B_V_dout,
        sync_nent => IL_L6PHID_neg2S_3_B_start,
        nent_o    => IL_L6PHID_neg2S_3_B_AV_dout_nent
      );

    IL_L6PHID_neg2S_3_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHID_neg2S_3_B_wea,
        addra     => IL_L6PHID_neg2S_3_B_writeaddr,
        dina      => IL_L6PHID_neg2S_3_B_din,
        wea_out       => IL_L6PHID_neg2S_3_B_wea_delay,
        addra_out     => IL_L6PHID_neg2S_3_B_writeaddr_delay,
        dina_out      => IL_L6PHID_neg2S_3_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHID_neg2S_3_B_start
      );

    IL_L6PHIA_neg2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIA_neg2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIA_neg2S_4_A_wea_delay,
        addra     => IL_L6PHIA_neg2S_4_A_writeaddr_delay,
        dina      => IL_L6PHIA_neg2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIA_neg2S_4_A_V_readaddr,
        doutb     => IL_L6PHIA_neg2S_4_A_V_dout,
        sync_nent => IL_L6PHIA_neg2S_4_A_start,
        nent_o    => IL_L6PHIA_neg2S_4_A_AV_dout_nent
      );

    IL_L6PHIA_neg2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIA_neg2S_4_A_wea,
        addra     => IL_L6PHIA_neg2S_4_A_writeaddr,
        dina      => IL_L6PHIA_neg2S_4_A_din,
        wea_out       => IL_L6PHIA_neg2S_4_A_wea_delay,
        addra_out     => IL_L6PHIA_neg2S_4_A_writeaddr_delay,
        dina_out      => IL_L6PHIA_neg2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIA_neg2S_4_A_start
      );

    IL_L6PHIB_neg2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIB_neg2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIB_neg2S_4_A_wea_delay,
        addra     => IL_L6PHIB_neg2S_4_A_writeaddr_delay,
        dina      => IL_L6PHIB_neg2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIB_neg2S_4_A_V_readaddr,
        doutb     => IL_L6PHIB_neg2S_4_A_V_dout,
        sync_nent => IL_L6PHIB_neg2S_4_A_start,
        nent_o    => IL_L6PHIB_neg2S_4_A_AV_dout_nent
      );

    IL_L6PHIB_neg2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIB_neg2S_4_A_wea,
        addra     => IL_L6PHIB_neg2S_4_A_writeaddr,
        dina      => IL_L6PHIB_neg2S_4_A_din,
        wea_out       => IL_L6PHIB_neg2S_4_A_wea_delay,
        addra_out     => IL_L6PHIB_neg2S_4_A_writeaddr_delay,
        dina_out      => IL_L6PHIB_neg2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_L6PHIB_neg2S_4_A_start
      );

    IL_L6PHIB_neg2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIB_neg2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIB_neg2S_4_B_wea_delay,
        addra     => IL_L6PHIB_neg2S_4_B_writeaddr_delay,
        dina      => IL_L6PHIB_neg2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIB_neg2S_4_B_V_readaddr,
        doutb     => IL_L6PHIB_neg2S_4_B_V_dout,
        sync_nent => IL_L6PHIB_neg2S_4_B_start,
        nent_o    => IL_L6PHIB_neg2S_4_B_AV_dout_nent
      );

    IL_L6PHIB_neg2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIB_neg2S_4_B_wea,
        addra     => IL_L6PHIB_neg2S_4_B_writeaddr,
        dina      => IL_L6PHIB_neg2S_4_B_din,
        wea_out       => IL_L6PHIB_neg2S_4_B_wea_delay,
        addra_out     => IL_L6PHIB_neg2S_4_B_writeaddr_delay,
        dina_out      => IL_L6PHIB_neg2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHIB_neg2S_4_B_start
      );

    IL_L6PHIC_neg2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHIC_neg2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHIC_neg2S_4_B_wea_delay,
        addra     => IL_L6PHIC_neg2S_4_B_writeaddr_delay,
        dina      => IL_L6PHIC_neg2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHIC_neg2S_4_B_V_readaddr,
        doutb     => IL_L6PHIC_neg2S_4_B_V_dout,
        sync_nent => IL_L6PHIC_neg2S_4_B_start,
        nent_o    => IL_L6PHIC_neg2S_4_B_AV_dout_nent
      );

    IL_L6PHIC_neg2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHIC_neg2S_4_B_wea,
        addra     => IL_L6PHIC_neg2S_4_B_writeaddr,
        dina      => IL_L6PHIC_neg2S_4_B_din,
        wea_out       => IL_L6PHIC_neg2S_4_B_wea_delay,
        addra_out     => IL_L6PHIC_neg2S_4_B_writeaddr_delay,
        dina_out      => IL_L6PHIC_neg2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHIC_neg2S_4_B_start
      );

    IL_L6PHID_neg2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_L6PHID_neg2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_L6PHID_neg2S_4_B_wea_delay,
        addra     => IL_L6PHID_neg2S_4_B_writeaddr_delay,
        dina      => IL_L6PHID_neg2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_L6PHID_neg2S_4_B_V_readaddr,
        doutb     => IL_L6PHID_neg2S_4_B_V_dout,
        sync_nent => IL_L6PHID_neg2S_4_B_start,
        nent_o    => IL_L6PHID_neg2S_4_B_AV_dout_nent
      );

    IL_L6PHID_neg2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_L6PHID_neg2S_4_B_wea,
        addra     => IL_L6PHID_neg2S_4_B_writeaddr,
        dina      => IL_L6PHID_neg2S_4_B_din,
        wea_out       => IL_L6PHID_neg2S_4_B_wea_delay,
        addra_out     => IL_L6PHID_neg2S_4_B_writeaddr_delay,
        dina_out      => IL_L6PHID_neg2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_L6PHID_neg2S_4_B_start
      );

    IL_D3PHIA_neg2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIA_neg2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIA_neg2S_4_A_wea_delay,
        addra     => IL_D3PHIA_neg2S_4_A_writeaddr_delay,
        dina      => IL_D3PHIA_neg2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIA_neg2S_4_A_V_readaddr,
        doutb     => IL_D3PHIA_neg2S_4_A_V_dout,
        sync_nent => IL_D3PHIA_neg2S_4_A_start,
        nent_o    => IL_D3PHIA_neg2S_4_A_AV_dout_nent
      );

    IL_D3PHIA_neg2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIA_neg2S_4_A_wea,
        addra     => IL_D3PHIA_neg2S_4_A_writeaddr,
        dina      => IL_D3PHIA_neg2S_4_A_din,
        wea_out       => IL_D3PHIA_neg2S_4_A_wea_delay,
        addra_out     => IL_D3PHIA_neg2S_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIA_neg2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIA_neg2S_4_A_start
      );

    IL_D3PHIB_neg2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_neg2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_neg2S_4_A_wea_delay,
        addra     => IL_D3PHIB_neg2S_4_A_writeaddr_delay,
        dina      => IL_D3PHIB_neg2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_neg2S_4_A_V_readaddr,
        doutb     => IL_D3PHIB_neg2S_4_A_V_dout,
        sync_nent => IL_D3PHIB_neg2S_4_A_start,
        nent_o    => IL_D3PHIB_neg2S_4_A_AV_dout_nent
      );

    IL_D3PHIB_neg2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_neg2S_4_A_wea,
        addra     => IL_D3PHIB_neg2S_4_A_writeaddr,
        dina      => IL_D3PHIB_neg2S_4_A_din,
        wea_out       => IL_D3PHIB_neg2S_4_A_wea_delay,
        addra_out     => IL_D3PHIB_neg2S_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIB_neg2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_neg2S_4_A_start
      );

    IL_D3PHIB_neg2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIB_neg2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIB_neg2S_4_B_wea_delay,
        addra     => IL_D3PHIB_neg2S_4_B_writeaddr_delay,
        dina      => IL_D3PHIB_neg2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIB_neg2S_4_B_V_readaddr,
        doutb     => IL_D3PHIB_neg2S_4_B_V_dout,
        sync_nent => IL_D3PHIB_neg2S_4_B_start,
        nent_o    => IL_D3PHIB_neg2S_4_B_AV_dout_nent
      );

    IL_D3PHIB_neg2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIB_neg2S_4_B_wea,
        addra     => IL_D3PHIB_neg2S_4_B_writeaddr,
        dina      => IL_D3PHIB_neg2S_4_B_din,
        wea_out       => IL_D3PHIB_neg2S_4_B_wea_delay,
        addra_out     => IL_D3PHIB_neg2S_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIB_neg2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIB_neg2S_4_B_start
      );

    IL_D3PHIC_neg2S_4_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_neg2S_4_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_neg2S_4_A_wea_delay,
        addra     => IL_D3PHIC_neg2S_4_A_writeaddr_delay,
        dina      => IL_D3PHIC_neg2S_4_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_neg2S_4_A_V_readaddr,
        doutb     => IL_D3PHIC_neg2S_4_A_V_dout,
        sync_nent => IL_D3PHIC_neg2S_4_A_start,
        nent_o    => IL_D3PHIC_neg2S_4_A_AV_dout_nent
      );

    IL_D3PHIC_neg2S_4_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_neg2S_4_A_wea,
        addra     => IL_D3PHIC_neg2S_4_A_writeaddr,
        dina      => IL_D3PHIC_neg2S_4_A_din,
        wea_out       => IL_D3PHIC_neg2S_4_A_wea_delay,
        addra_out     => IL_D3PHIC_neg2S_4_A_writeaddr_delay,
        dina_out      => IL_D3PHIC_neg2S_4_A_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_neg2S_4_A_start
      );

    IL_D3PHIC_neg2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHIC_neg2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHIC_neg2S_4_B_wea_delay,
        addra     => IL_D3PHIC_neg2S_4_B_writeaddr_delay,
        dina      => IL_D3PHIC_neg2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHIC_neg2S_4_B_V_readaddr,
        doutb     => IL_D3PHIC_neg2S_4_B_V_dout,
        sync_nent => IL_D3PHIC_neg2S_4_B_start,
        nent_o    => IL_D3PHIC_neg2S_4_B_AV_dout_nent
      );

    IL_D3PHIC_neg2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHIC_neg2S_4_B_wea,
        addra     => IL_D3PHIC_neg2S_4_B_writeaddr,
        dina      => IL_D3PHIC_neg2S_4_B_din,
        wea_out       => IL_D3PHIC_neg2S_4_B_wea_delay,
        addra_out     => IL_D3PHIC_neg2S_4_B_writeaddr_delay,
        dina_out      => IL_D3PHIC_neg2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHIC_neg2S_4_B_start
      );

    IL_D3PHID_neg2S_4_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D3PHID_neg2S_4_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D3PHID_neg2S_4_B_wea_delay,
        addra     => IL_D3PHID_neg2S_4_B_writeaddr_delay,
        dina      => IL_D3PHID_neg2S_4_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D3PHID_neg2S_4_B_V_readaddr,
        doutb     => IL_D3PHID_neg2S_4_B_V_dout,
        sync_nent => IL_D3PHID_neg2S_4_B_start,
        nent_o    => IL_D3PHID_neg2S_4_B_AV_dout_nent
      );

    IL_D3PHID_neg2S_4_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D3PHID_neg2S_4_B_wea,
        addra     => IL_D3PHID_neg2S_4_B_writeaddr,
        dina      => IL_D3PHID_neg2S_4_B_din,
        wea_out       => IL_D3PHID_neg2S_4_B_wea_delay,
        addra_out     => IL_D3PHID_neg2S_4_B_writeaddr_delay,
        dina_out      => IL_D3PHID_neg2S_4_B_din_delay,
        done       => IR_done,
        start      => IL_D3PHID_neg2S_4_B_start
      );

    IL_D1PHIA_neg2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIA_neg2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIA_neg2S_5_A_wea_delay,
        addra     => IL_D1PHIA_neg2S_5_A_writeaddr_delay,
        dina      => IL_D1PHIA_neg2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIA_neg2S_5_A_V_readaddr,
        doutb     => IL_D1PHIA_neg2S_5_A_V_dout,
        sync_nent => IL_D1PHIA_neg2S_5_A_start,
        nent_o    => IL_D1PHIA_neg2S_5_A_AV_dout_nent
      );

    IL_D1PHIA_neg2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIA_neg2S_5_A_wea,
        addra     => IL_D1PHIA_neg2S_5_A_writeaddr,
        dina      => IL_D1PHIA_neg2S_5_A_din,
        wea_out       => IL_D1PHIA_neg2S_5_A_wea_delay,
        addra_out     => IL_D1PHIA_neg2S_5_A_writeaddr_delay,
        dina_out      => IL_D1PHIA_neg2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIA_neg2S_5_A_start
      );

    IL_D1PHIB_neg2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_neg2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_neg2S_5_A_wea_delay,
        addra     => IL_D1PHIB_neg2S_5_A_writeaddr_delay,
        dina      => IL_D1PHIB_neg2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_neg2S_5_A_V_readaddr,
        doutb     => IL_D1PHIB_neg2S_5_A_V_dout,
        sync_nent => IL_D1PHIB_neg2S_5_A_start,
        nent_o    => IL_D1PHIB_neg2S_5_A_AV_dout_nent
      );

    IL_D1PHIB_neg2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_neg2S_5_A_wea,
        addra     => IL_D1PHIB_neg2S_5_A_writeaddr,
        dina      => IL_D1PHIB_neg2S_5_A_din,
        wea_out       => IL_D1PHIB_neg2S_5_A_wea_delay,
        addra_out     => IL_D1PHIB_neg2S_5_A_writeaddr_delay,
        dina_out      => IL_D1PHIB_neg2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_neg2S_5_A_start
      );

    IL_D1PHIB_neg2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIB_neg2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIB_neg2S_5_B_wea_delay,
        addra     => IL_D1PHIB_neg2S_5_B_writeaddr_delay,
        dina      => IL_D1PHIB_neg2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIB_neg2S_5_B_V_readaddr,
        doutb     => IL_D1PHIB_neg2S_5_B_V_dout,
        sync_nent => IL_D1PHIB_neg2S_5_B_start,
        nent_o    => IL_D1PHIB_neg2S_5_B_AV_dout_nent
      );

    IL_D1PHIB_neg2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIB_neg2S_5_B_wea,
        addra     => IL_D1PHIB_neg2S_5_B_writeaddr,
        dina      => IL_D1PHIB_neg2S_5_B_din,
        wea_out       => IL_D1PHIB_neg2S_5_B_wea_delay,
        addra_out     => IL_D1PHIB_neg2S_5_B_writeaddr_delay,
        dina_out      => IL_D1PHIB_neg2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIB_neg2S_5_B_start
      );

    IL_D1PHIC_neg2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_neg2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_neg2S_5_A_wea_delay,
        addra     => IL_D1PHIC_neg2S_5_A_writeaddr_delay,
        dina      => IL_D1PHIC_neg2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_neg2S_5_A_V_readaddr,
        doutb     => IL_D1PHIC_neg2S_5_A_V_dout,
        sync_nent => IL_D1PHIC_neg2S_5_A_start,
        nent_o    => IL_D1PHIC_neg2S_5_A_AV_dout_nent
      );

    IL_D1PHIC_neg2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_neg2S_5_A_wea,
        addra     => IL_D1PHIC_neg2S_5_A_writeaddr,
        dina      => IL_D1PHIC_neg2S_5_A_din,
        wea_out       => IL_D1PHIC_neg2S_5_A_wea_delay,
        addra_out     => IL_D1PHIC_neg2S_5_A_writeaddr_delay,
        dina_out      => IL_D1PHIC_neg2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_neg2S_5_A_start
      );

    IL_D1PHIC_neg2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHIC_neg2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHIC_neg2S_5_B_wea_delay,
        addra     => IL_D1PHIC_neg2S_5_B_writeaddr_delay,
        dina      => IL_D1PHIC_neg2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHIC_neg2S_5_B_V_readaddr,
        doutb     => IL_D1PHIC_neg2S_5_B_V_dout,
        sync_nent => IL_D1PHIC_neg2S_5_B_start,
        nent_o    => IL_D1PHIC_neg2S_5_B_AV_dout_nent
      );

    IL_D1PHIC_neg2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHIC_neg2S_5_B_wea,
        addra     => IL_D1PHIC_neg2S_5_B_writeaddr,
        dina      => IL_D1PHIC_neg2S_5_B_din,
        wea_out       => IL_D1PHIC_neg2S_5_B_wea_delay,
        addra_out     => IL_D1PHIC_neg2S_5_B_writeaddr_delay,
        dina_out      => IL_D1PHIC_neg2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHIC_neg2S_5_B_start
      );

    IL_D1PHID_neg2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D1PHID_neg2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D1PHID_neg2S_5_B_wea_delay,
        addra     => IL_D1PHID_neg2S_5_B_writeaddr_delay,
        dina      => IL_D1PHID_neg2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D1PHID_neg2S_5_B_V_readaddr,
        doutb     => IL_D1PHID_neg2S_5_B_V_dout,
        sync_nent => IL_D1PHID_neg2S_5_B_start,
        nent_o    => IL_D1PHID_neg2S_5_B_AV_dout_nent
      );

    IL_D1PHID_neg2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D1PHID_neg2S_5_B_wea,
        addra     => IL_D1PHID_neg2S_5_B_writeaddr,
        dina      => IL_D1PHID_neg2S_5_B_din,
        wea_out       => IL_D1PHID_neg2S_5_B_wea_delay,
        addra_out     => IL_D1PHID_neg2S_5_B_writeaddr_delay,
        dina_out      => IL_D1PHID_neg2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D1PHID_neg2S_5_B_start
      );

    IL_D4PHIA_neg2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIA_neg2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIA_neg2S_5_A_wea_delay,
        addra     => IL_D4PHIA_neg2S_5_A_writeaddr_delay,
        dina      => IL_D4PHIA_neg2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIA_neg2S_5_A_V_readaddr,
        doutb     => IL_D4PHIA_neg2S_5_A_V_dout,
        sync_nent => IL_D4PHIA_neg2S_5_A_start,
        nent_o    => IL_D4PHIA_neg2S_5_A_AV_dout_nent
      );

    IL_D4PHIA_neg2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIA_neg2S_5_A_wea,
        addra     => IL_D4PHIA_neg2S_5_A_writeaddr,
        dina      => IL_D4PHIA_neg2S_5_A_din,
        wea_out       => IL_D4PHIA_neg2S_5_A_wea_delay,
        addra_out     => IL_D4PHIA_neg2S_5_A_writeaddr_delay,
        dina_out      => IL_D4PHIA_neg2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIA_neg2S_5_A_start
      );

    IL_D4PHIB_neg2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_neg2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_neg2S_5_A_wea_delay,
        addra     => IL_D4PHIB_neg2S_5_A_writeaddr_delay,
        dina      => IL_D4PHIB_neg2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_neg2S_5_A_V_readaddr,
        doutb     => IL_D4PHIB_neg2S_5_A_V_dout,
        sync_nent => IL_D4PHIB_neg2S_5_A_start,
        nent_o    => IL_D4PHIB_neg2S_5_A_AV_dout_nent
      );

    IL_D4PHIB_neg2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_neg2S_5_A_wea,
        addra     => IL_D4PHIB_neg2S_5_A_writeaddr,
        dina      => IL_D4PHIB_neg2S_5_A_din,
        wea_out       => IL_D4PHIB_neg2S_5_A_wea_delay,
        addra_out     => IL_D4PHIB_neg2S_5_A_writeaddr_delay,
        dina_out      => IL_D4PHIB_neg2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_neg2S_5_A_start
      );

    IL_D4PHIB_neg2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIB_neg2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIB_neg2S_5_B_wea_delay,
        addra     => IL_D4PHIB_neg2S_5_B_writeaddr_delay,
        dina      => IL_D4PHIB_neg2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIB_neg2S_5_B_V_readaddr,
        doutb     => IL_D4PHIB_neg2S_5_B_V_dout,
        sync_nent => IL_D4PHIB_neg2S_5_B_start,
        nent_o    => IL_D4PHIB_neg2S_5_B_AV_dout_nent
      );

    IL_D4PHIB_neg2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIB_neg2S_5_B_wea,
        addra     => IL_D4PHIB_neg2S_5_B_writeaddr,
        dina      => IL_D4PHIB_neg2S_5_B_din,
        wea_out       => IL_D4PHIB_neg2S_5_B_wea_delay,
        addra_out     => IL_D4PHIB_neg2S_5_B_writeaddr_delay,
        dina_out      => IL_D4PHIB_neg2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIB_neg2S_5_B_start
      );

    IL_D4PHIC_neg2S_5_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_neg2S_5_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_neg2S_5_A_wea_delay,
        addra     => IL_D4PHIC_neg2S_5_A_writeaddr_delay,
        dina      => IL_D4PHIC_neg2S_5_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_neg2S_5_A_V_readaddr,
        doutb     => IL_D4PHIC_neg2S_5_A_V_dout,
        sync_nent => IL_D4PHIC_neg2S_5_A_start,
        nent_o    => IL_D4PHIC_neg2S_5_A_AV_dout_nent
      );

    IL_D4PHIC_neg2S_5_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_neg2S_5_A_wea,
        addra     => IL_D4PHIC_neg2S_5_A_writeaddr,
        dina      => IL_D4PHIC_neg2S_5_A_din,
        wea_out       => IL_D4PHIC_neg2S_5_A_wea_delay,
        addra_out     => IL_D4PHIC_neg2S_5_A_writeaddr_delay,
        dina_out      => IL_D4PHIC_neg2S_5_A_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_neg2S_5_A_start
      );

    IL_D4PHIC_neg2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHIC_neg2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHIC_neg2S_5_B_wea_delay,
        addra     => IL_D4PHIC_neg2S_5_B_writeaddr_delay,
        dina      => IL_D4PHIC_neg2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHIC_neg2S_5_B_V_readaddr,
        doutb     => IL_D4PHIC_neg2S_5_B_V_dout,
        sync_nent => IL_D4PHIC_neg2S_5_B_start,
        nent_o    => IL_D4PHIC_neg2S_5_B_AV_dout_nent
      );

    IL_D4PHIC_neg2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHIC_neg2S_5_B_wea,
        addra     => IL_D4PHIC_neg2S_5_B_writeaddr,
        dina      => IL_D4PHIC_neg2S_5_B_din,
        wea_out       => IL_D4PHIC_neg2S_5_B_wea_delay,
        addra_out     => IL_D4PHIC_neg2S_5_B_writeaddr_delay,
        dina_out      => IL_D4PHIC_neg2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHIC_neg2S_5_B_start
      );

    IL_D4PHID_neg2S_5_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D4PHID_neg2S_5_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D4PHID_neg2S_5_B_wea_delay,
        addra     => IL_D4PHID_neg2S_5_B_writeaddr_delay,
        dina      => IL_D4PHID_neg2S_5_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D4PHID_neg2S_5_B_V_readaddr,
        doutb     => IL_D4PHID_neg2S_5_B_V_dout,
        sync_nent => IL_D4PHID_neg2S_5_B_start,
        nent_o    => IL_D4PHID_neg2S_5_B_AV_dout_nent
      );

    IL_D4PHID_neg2S_5_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D4PHID_neg2S_5_B_wea,
        addra     => IL_D4PHID_neg2S_5_B_writeaddr,
        dina      => IL_D4PHID_neg2S_5_B_din,
        wea_out       => IL_D4PHID_neg2S_5_B_wea_delay,
        addra_out     => IL_D4PHID_neg2S_5_B_writeaddr_delay,
        dina_out      => IL_D4PHID_neg2S_5_B_din_delay,
        done       => IR_done,
        start      => IL_D4PHID_neg2S_5_B_start
      );

    IL_D2PHIA_neg2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIA_neg2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIA_neg2S_6_A_wea_delay,
        addra     => IL_D2PHIA_neg2S_6_A_writeaddr_delay,
        dina      => IL_D2PHIA_neg2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIA_neg2S_6_A_V_readaddr,
        doutb     => IL_D2PHIA_neg2S_6_A_V_dout,
        sync_nent => IL_D2PHIA_neg2S_6_A_start,
        nent_o    => IL_D2PHIA_neg2S_6_A_AV_dout_nent
      );

    IL_D2PHIA_neg2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIA_neg2S_6_A_wea,
        addra     => IL_D2PHIA_neg2S_6_A_writeaddr,
        dina      => IL_D2PHIA_neg2S_6_A_din,
        wea_out       => IL_D2PHIA_neg2S_6_A_wea_delay,
        addra_out     => IL_D2PHIA_neg2S_6_A_writeaddr_delay,
        dina_out      => IL_D2PHIA_neg2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIA_neg2S_6_A_start
      );

    IL_D2PHIB_neg2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_neg2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_neg2S_6_A_wea_delay,
        addra     => IL_D2PHIB_neg2S_6_A_writeaddr_delay,
        dina      => IL_D2PHIB_neg2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_neg2S_6_A_V_readaddr,
        doutb     => IL_D2PHIB_neg2S_6_A_V_dout,
        sync_nent => IL_D2PHIB_neg2S_6_A_start,
        nent_o    => IL_D2PHIB_neg2S_6_A_AV_dout_nent
      );

    IL_D2PHIB_neg2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_neg2S_6_A_wea,
        addra     => IL_D2PHIB_neg2S_6_A_writeaddr,
        dina      => IL_D2PHIB_neg2S_6_A_din,
        wea_out       => IL_D2PHIB_neg2S_6_A_wea_delay,
        addra_out     => IL_D2PHIB_neg2S_6_A_writeaddr_delay,
        dina_out      => IL_D2PHIB_neg2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_neg2S_6_A_start
      );

    IL_D2PHIB_neg2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIB_neg2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIB_neg2S_6_B_wea_delay,
        addra     => IL_D2PHIB_neg2S_6_B_writeaddr_delay,
        dina      => IL_D2PHIB_neg2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIB_neg2S_6_B_V_readaddr,
        doutb     => IL_D2PHIB_neg2S_6_B_V_dout,
        sync_nent => IL_D2PHIB_neg2S_6_B_start,
        nent_o    => IL_D2PHIB_neg2S_6_B_AV_dout_nent
      );

    IL_D2PHIB_neg2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIB_neg2S_6_B_wea,
        addra     => IL_D2PHIB_neg2S_6_B_writeaddr,
        dina      => IL_D2PHIB_neg2S_6_B_din,
        wea_out       => IL_D2PHIB_neg2S_6_B_wea_delay,
        addra_out     => IL_D2PHIB_neg2S_6_B_writeaddr_delay,
        dina_out      => IL_D2PHIB_neg2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIB_neg2S_6_B_start
      );

    IL_D2PHIC_neg2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_neg2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_neg2S_6_A_wea_delay,
        addra     => IL_D2PHIC_neg2S_6_A_writeaddr_delay,
        dina      => IL_D2PHIC_neg2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_neg2S_6_A_V_readaddr,
        doutb     => IL_D2PHIC_neg2S_6_A_V_dout,
        sync_nent => IL_D2PHIC_neg2S_6_A_start,
        nent_o    => IL_D2PHIC_neg2S_6_A_AV_dout_nent
      );

    IL_D2PHIC_neg2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_neg2S_6_A_wea,
        addra     => IL_D2PHIC_neg2S_6_A_writeaddr,
        dina      => IL_D2PHIC_neg2S_6_A_din,
        wea_out       => IL_D2PHIC_neg2S_6_A_wea_delay,
        addra_out     => IL_D2PHIC_neg2S_6_A_writeaddr_delay,
        dina_out      => IL_D2PHIC_neg2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_neg2S_6_A_start
      );

    IL_D2PHIC_neg2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHIC_neg2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHIC_neg2S_6_B_wea_delay,
        addra     => IL_D2PHIC_neg2S_6_B_writeaddr_delay,
        dina      => IL_D2PHIC_neg2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHIC_neg2S_6_B_V_readaddr,
        doutb     => IL_D2PHIC_neg2S_6_B_V_dout,
        sync_nent => IL_D2PHIC_neg2S_6_B_start,
        nent_o    => IL_D2PHIC_neg2S_6_B_AV_dout_nent
      );

    IL_D2PHIC_neg2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHIC_neg2S_6_B_wea,
        addra     => IL_D2PHIC_neg2S_6_B_writeaddr,
        dina      => IL_D2PHIC_neg2S_6_B_din,
        wea_out       => IL_D2PHIC_neg2S_6_B_wea_delay,
        addra_out     => IL_D2PHIC_neg2S_6_B_writeaddr_delay,
        dina_out      => IL_D2PHIC_neg2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHIC_neg2S_6_B_start
      );

    IL_D2PHID_neg2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D2PHID_neg2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D2PHID_neg2S_6_B_wea_delay,
        addra     => IL_D2PHID_neg2S_6_B_writeaddr_delay,
        dina      => IL_D2PHID_neg2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D2PHID_neg2S_6_B_V_readaddr,
        doutb     => IL_D2PHID_neg2S_6_B_V_dout,
        sync_nent => IL_D2PHID_neg2S_6_B_start,
        nent_o    => IL_D2PHID_neg2S_6_B_AV_dout_nent
      );

    IL_D2PHID_neg2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D2PHID_neg2S_6_B_wea,
        addra     => IL_D2PHID_neg2S_6_B_writeaddr,
        dina      => IL_D2PHID_neg2S_6_B_din,
        wea_out       => IL_D2PHID_neg2S_6_B_wea_delay,
        addra_out     => IL_D2PHID_neg2S_6_B_writeaddr_delay,
        dina_out      => IL_D2PHID_neg2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D2PHID_neg2S_6_B_start
      );

    IL_D5PHIA_neg2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIA_neg2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIA_neg2S_6_A_wea_delay,
        addra     => IL_D5PHIA_neg2S_6_A_writeaddr_delay,
        dina      => IL_D5PHIA_neg2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIA_neg2S_6_A_V_readaddr,
        doutb     => IL_D5PHIA_neg2S_6_A_V_dout,
        sync_nent => IL_D5PHIA_neg2S_6_A_start,
        nent_o    => IL_D5PHIA_neg2S_6_A_AV_dout_nent
      );

    IL_D5PHIA_neg2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIA_neg2S_6_A_wea,
        addra     => IL_D5PHIA_neg2S_6_A_writeaddr,
        dina      => IL_D5PHIA_neg2S_6_A_din,
        wea_out       => IL_D5PHIA_neg2S_6_A_wea_delay,
        addra_out     => IL_D5PHIA_neg2S_6_A_writeaddr_delay,
        dina_out      => IL_D5PHIA_neg2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIA_neg2S_6_A_start
      );

    IL_D5PHIB_neg2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_neg2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_neg2S_6_A_wea_delay,
        addra     => IL_D5PHIB_neg2S_6_A_writeaddr_delay,
        dina      => IL_D5PHIB_neg2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_neg2S_6_A_V_readaddr,
        doutb     => IL_D5PHIB_neg2S_6_A_V_dout,
        sync_nent => IL_D5PHIB_neg2S_6_A_start,
        nent_o    => IL_D5PHIB_neg2S_6_A_AV_dout_nent
      );

    IL_D5PHIB_neg2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_neg2S_6_A_wea,
        addra     => IL_D5PHIB_neg2S_6_A_writeaddr,
        dina      => IL_D5PHIB_neg2S_6_A_din,
        wea_out       => IL_D5PHIB_neg2S_6_A_wea_delay,
        addra_out     => IL_D5PHIB_neg2S_6_A_writeaddr_delay,
        dina_out      => IL_D5PHIB_neg2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_neg2S_6_A_start
      );

    IL_D5PHIB_neg2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIB_neg2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIB_neg2S_6_B_wea_delay,
        addra     => IL_D5PHIB_neg2S_6_B_writeaddr_delay,
        dina      => IL_D5PHIB_neg2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIB_neg2S_6_B_V_readaddr,
        doutb     => IL_D5PHIB_neg2S_6_B_V_dout,
        sync_nent => IL_D5PHIB_neg2S_6_B_start,
        nent_o    => IL_D5PHIB_neg2S_6_B_AV_dout_nent
      );

    IL_D5PHIB_neg2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIB_neg2S_6_B_wea,
        addra     => IL_D5PHIB_neg2S_6_B_writeaddr,
        dina      => IL_D5PHIB_neg2S_6_B_din,
        wea_out       => IL_D5PHIB_neg2S_6_B_wea_delay,
        addra_out     => IL_D5PHIB_neg2S_6_B_writeaddr_delay,
        dina_out      => IL_D5PHIB_neg2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIB_neg2S_6_B_start
      );

    IL_D5PHIC_neg2S_6_A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_neg2S_6_A"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_neg2S_6_A_wea_delay,
        addra     => IL_D5PHIC_neg2S_6_A_writeaddr_delay,
        dina      => IL_D5PHIC_neg2S_6_A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_neg2S_6_A_V_readaddr,
        doutb     => IL_D5PHIC_neg2S_6_A_V_dout,
        sync_nent => IL_D5PHIC_neg2S_6_A_start,
        nent_o    => IL_D5PHIC_neg2S_6_A_AV_dout_nent
      );

    IL_D5PHIC_neg2S_6_A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_neg2S_6_A_wea,
        addra     => IL_D5PHIC_neg2S_6_A_writeaddr,
        dina      => IL_D5PHIC_neg2S_6_A_din,
        wea_out       => IL_D5PHIC_neg2S_6_A_wea_delay,
        addra_out     => IL_D5PHIC_neg2S_6_A_writeaddr_delay,
        dina_out      => IL_D5PHIC_neg2S_6_A_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_neg2S_6_A_start
      );

    IL_D5PHIC_neg2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHIC_neg2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHIC_neg2S_6_B_wea_delay,
        addra     => IL_D5PHIC_neg2S_6_B_writeaddr_delay,
        dina      => IL_D5PHIC_neg2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHIC_neg2S_6_B_V_readaddr,
        doutb     => IL_D5PHIC_neg2S_6_B_V_dout,
        sync_nent => IL_D5PHIC_neg2S_6_B_start,
        nent_o    => IL_D5PHIC_neg2S_6_B_AV_dout_nent
      );

    IL_D5PHIC_neg2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHIC_neg2S_6_B_wea,
        addra     => IL_D5PHIC_neg2S_6_B_writeaddr,
        dina      => IL_D5PHIC_neg2S_6_B_din,
        wea_out       => IL_D5PHIC_neg2S_6_B_wea_delay,
        addra_out     => IL_D5PHIC_neg2S_6_B_writeaddr_delay,
        dina_out      => IL_D5PHIC_neg2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHIC_neg2S_6_B_start
      );

    IL_D5PHID_neg2S_6_B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "IL_D5PHID_neg2S_6_B"
      )
      port map (
        clka      => clk,
        wea       => IL_D5PHID_neg2S_6_B_wea_delay,
        addra     => IL_D5PHID_neg2S_6_B_writeaddr_delay,
        dina      => IL_D5PHID_neg2S_6_B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => IL_D5PHID_neg2S_6_B_V_readaddr,
        doutb     => IL_D5PHID_neg2S_6_B_V_dout,
        sync_nent => IL_D5PHID_neg2S_6_B_start,
        nent_o    => IL_D5PHID_neg2S_6_B_AV_dout_nent
      );

    IL_D5PHID_neg2S_6_B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => IL_D5PHID_neg2S_6_B_wea,
        addra     => IL_D5PHID_neg2S_6_B_writeaddr,
        dina      => IL_D5PHID_neg2S_6_B_din,
        wea_out       => IL_D5PHID_neg2S_6_B_wea_delay,
        addra_out     => IL_D5PHID_neg2S_6_B_writeaddr_delay,
        dina_out      => IL_D5PHID_neg2S_6_B_din_delay,
        done       => IR_done,
        start      => IL_D5PHID_neg2S_6_B_start
      );

    AS_L1PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHIAn1_bx,
        bx_vld => AS_L1PHIAn1_bx_vld
      );

--    STREAM_AS_L1PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHIAn1_bx,
--        bx_in_vld => AS_L1PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHIAn1_stream_V_dout,
--        din0=>AS_L1PHIAn1_V_dout,
--        din1=>AS_L1PHIAn1_V_dout,
--        din2=>AS_L1PHIAn1_V_dout,
--        din3=>AS_L1PHIAn1_V_dout,
--        nent0=>AS_L1PHIAn1_AV_dout_nent,
--        nent1=>AS_L1PHIAn1_AV_dout_nent,
--        nent2=>AS_L1PHIAn1_AV_dout_nent,
--        nent3=>AS_L1PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHIAn1_V_readaddr
--      );

    AS_L1PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIAn1_wea_delay,
        addra     => AS_L1PHIAn1_writeaddr_delay,
        dina      => AS_L1PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIAn1_V_readaddr,
        doutb     => AS_L1PHIAn1_V_dout,
        sync_nent => AS_L1PHIAn1_start,
        nent_o    => AS_L1PHIAn1_AV_dout_nent
      );

    AS_L1PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIAn1_wea,
        addra     => AS_L1PHIAn1_writeaddr,
        dina      => AS_L1PHIAn1_din,
        wea_out       => AS_L1PHIAn1_wea_delay,
        addra_out     => AS_L1PHIAn1_writeaddr_delay,
        dina_out      => AS_L1PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIAn1_start
      );

    AS_L1PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHIBn1_bx,
        bx_vld => AS_L1PHIBn1_bx_vld
      );

--    STREAM_AS_L1PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHIBn1_bx,
--        bx_in_vld => AS_L1PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHIBn1_stream_V_dout,
--        din0=>AS_L1PHIBn1_V_dout,
--        din1=>AS_L1PHIBn1_V_dout,
--        din2=>AS_L1PHIBn1_V_dout,
--        din3=>AS_L1PHIBn1_V_dout,
--        nent0=>AS_L1PHIBn1_AV_dout_nent,
--        nent1=>AS_L1PHIBn1_AV_dout_nent,
--        nent2=>AS_L1PHIBn1_AV_dout_nent,
--        nent3=>AS_L1PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHIBn1_V_readaddr
--      );

    AS_L1PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIBn1_wea_delay,
        addra     => AS_L1PHIBn1_writeaddr_delay,
        dina      => AS_L1PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIBn1_V_readaddr,
        doutb     => AS_L1PHIBn1_V_dout,
        sync_nent => AS_L1PHIBn1_start,
        nent_o    => AS_L1PHIBn1_AV_dout_nent
      );

    AS_L1PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIBn1_wea,
        addra     => AS_L1PHIBn1_writeaddr,
        dina      => AS_L1PHIBn1_din,
        wea_out       => AS_L1PHIBn1_wea_delay,
        addra_out     => AS_L1PHIBn1_writeaddr_delay,
        dina_out      => AS_L1PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIBn1_start
      );

    AS_L1PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHICn1_bx,
        bx_vld => AS_L1PHICn1_bx_vld
      );

--    STREAM_AS_L1PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHICn1_bx,
--        bx_in_vld => AS_L1PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHICn1_stream_V_dout,
--        din0=>AS_L1PHICn1_V_dout,
--        din1=>AS_L1PHICn1_V_dout,
--        din2=>AS_L1PHICn1_V_dout,
--        din3=>AS_L1PHICn1_V_dout,
--        nent0=>AS_L1PHICn1_AV_dout_nent,
--        nent1=>AS_L1PHICn1_AV_dout_nent,
--        nent2=>AS_L1PHICn1_AV_dout_nent,
--        nent3=>AS_L1PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHICn1_V_readaddr
--      );

    AS_L1PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHICn1_wea_delay,
        addra     => AS_L1PHICn1_writeaddr_delay,
        dina      => AS_L1PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHICn1_V_readaddr,
        doutb     => AS_L1PHICn1_V_dout,
        sync_nent => AS_L1PHICn1_start,
        nent_o    => AS_L1PHICn1_AV_dout_nent
      );

    AS_L1PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHICn1_wea,
        addra     => AS_L1PHICn1_writeaddr,
        dina      => AS_L1PHICn1_din,
        wea_out       => AS_L1PHICn1_wea_delay,
        addra_out     => AS_L1PHICn1_writeaddr_delay,
        dina_out      => AS_L1PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHICn1_start
      );

    AS_L1PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHIDn1_bx,
        bx_vld => AS_L1PHIDn1_bx_vld
      );

--    STREAM_AS_L1PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHIDn1_bx,
--        bx_in_vld => AS_L1PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHIDn1_stream_V_dout,
--        din0=>AS_L1PHIDn1_V_dout,
--        din1=>AS_L1PHIDn1_V_dout,
--        din2=>AS_L1PHIDn1_V_dout,
--        din3=>AS_L1PHIDn1_V_dout,
--        nent0=>AS_L1PHIDn1_AV_dout_nent,
--        nent1=>AS_L1PHIDn1_AV_dout_nent,
--        nent2=>AS_L1PHIDn1_AV_dout_nent,
--        nent3=>AS_L1PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHIDn1_V_readaddr
--      );

    AS_L1PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIDn1_wea_delay,
        addra     => AS_L1PHIDn1_writeaddr_delay,
        dina      => AS_L1PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIDn1_V_readaddr,
        doutb     => AS_L1PHIDn1_V_dout,
        sync_nent => AS_L1PHIDn1_start,
        nent_o    => AS_L1PHIDn1_AV_dout_nent
      );

    AS_L1PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIDn1_wea,
        addra     => AS_L1PHIDn1_writeaddr,
        dina      => AS_L1PHIDn1_din,
        wea_out       => AS_L1PHIDn1_wea_delay,
        addra_out     => AS_L1PHIDn1_writeaddr_delay,
        dina_out      => AS_L1PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIDn1_start
      );

    AS_L1PHIEn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHIEn1_bx,
        bx_vld => AS_L1PHIEn1_bx_vld
      );

--    STREAM_AS_L1PHIEn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHIEn1_bx,
--        bx_in_vld => AS_L1PHIEn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHIEn1_stream_V_dout,
--        din0=>AS_L1PHIEn1_V_dout,
--        din1=>AS_L1PHIEn1_V_dout,
--        din2=>AS_L1PHIEn1_V_dout,
--        din3=>AS_L1PHIEn1_V_dout,
--        nent0=>AS_L1PHIEn1_AV_dout_nent,
--        nent1=>AS_L1PHIEn1_AV_dout_nent,
--        nent2=>AS_L1PHIEn1_AV_dout_nent,
--        nent3=>AS_L1PHIEn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHIEn1_V_readaddr
--      );

    AS_L1PHIEn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIEn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIEn1_wea_delay,
        addra     => AS_L1PHIEn1_writeaddr_delay,
        dina      => AS_L1PHIEn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIEn1_V_readaddr,
        doutb     => AS_L1PHIEn1_V_dout,
        sync_nent => AS_L1PHIEn1_start,
        nent_o    => AS_L1PHIEn1_AV_dout_nent
      );

    AS_L1PHIEn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIEn1_wea,
        addra     => AS_L1PHIEn1_writeaddr,
        dina      => AS_L1PHIEn1_din,
        wea_out       => AS_L1PHIEn1_wea_delay,
        addra_out     => AS_L1PHIEn1_writeaddr_delay,
        dina_out      => AS_L1PHIEn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIEn1_start
      );

    AS_L1PHIFn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHIFn1_bx,
        bx_vld => AS_L1PHIFn1_bx_vld
      );

--    STREAM_AS_L1PHIFn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHIFn1_bx,
--        bx_in_vld => AS_L1PHIFn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHIFn1_stream_V_dout,
--        din0=>AS_L1PHIFn1_V_dout,
--        din1=>AS_L1PHIFn1_V_dout,
--        din2=>AS_L1PHIFn1_V_dout,
--        din3=>AS_L1PHIFn1_V_dout,
--        nent0=>AS_L1PHIFn1_AV_dout_nent,
--        nent1=>AS_L1PHIFn1_AV_dout_nent,
--        nent2=>AS_L1PHIFn1_AV_dout_nent,
--        nent3=>AS_L1PHIFn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHIFn1_V_readaddr
--      );

    AS_L1PHIFn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIFn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIFn1_wea_delay,
        addra     => AS_L1PHIFn1_writeaddr_delay,
        dina      => AS_L1PHIFn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIFn1_V_readaddr,
        doutb     => AS_L1PHIFn1_V_dout,
        sync_nent => AS_L1PHIFn1_start,
        nent_o    => AS_L1PHIFn1_AV_dout_nent
      );

    AS_L1PHIFn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIFn1_wea,
        addra     => AS_L1PHIFn1_writeaddr,
        dina      => AS_L1PHIFn1_din,
        wea_out       => AS_L1PHIFn1_wea_delay,
        addra_out     => AS_L1PHIFn1_writeaddr_delay,
        dina_out      => AS_L1PHIFn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIFn1_start
      );

    AS_L1PHIGn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHIGn1_bx,
        bx_vld => AS_L1PHIGn1_bx_vld
      );

--    STREAM_AS_L1PHIGn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHIGn1_bx,
--        bx_in_vld => AS_L1PHIGn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHIGn1_stream_V_dout,
--        din0=>AS_L1PHIGn1_V_dout,
--        din1=>AS_L1PHIGn1_V_dout,
--        din2=>AS_L1PHIGn1_V_dout,
--        din3=>AS_L1PHIGn1_V_dout,
--        nent0=>AS_L1PHIGn1_AV_dout_nent,
--        nent1=>AS_L1PHIGn1_AV_dout_nent,
--        nent2=>AS_L1PHIGn1_AV_dout_nent,
--        nent3=>AS_L1PHIGn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHIGn1_V_readaddr
--      );

    AS_L1PHIGn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIGn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIGn1_wea_delay,
        addra     => AS_L1PHIGn1_writeaddr_delay,
        dina      => AS_L1PHIGn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIGn1_V_readaddr,
        doutb     => AS_L1PHIGn1_V_dout,
        sync_nent => AS_L1PHIGn1_start,
        nent_o    => AS_L1PHIGn1_AV_dout_nent
      );

    AS_L1PHIGn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIGn1_wea,
        addra     => AS_L1PHIGn1_writeaddr,
        dina      => AS_L1PHIGn1_din,
        wea_out       => AS_L1PHIGn1_wea_delay,
        addra_out     => AS_L1PHIGn1_writeaddr_delay,
        dina_out      => AS_L1PHIGn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIGn1_start
      );

    AS_L1PHIHn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L1PHIHn1_bx,
        bx_vld => AS_L1PHIHn1_bx_vld
      );

--    STREAM_AS_L1PHIHn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L1PHIHn1_bx,
--        bx_in_vld => AS_L1PHIHn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L1PHIHn1_stream_V_dout,
--        din0=>AS_L1PHIHn1_V_dout,
--        din1=>AS_L1PHIHn1_V_dout,
--        din2=>AS_L1PHIHn1_V_dout,
--        din3=>AS_L1PHIHn1_V_dout,
--        nent0=>AS_L1PHIHn1_AV_dout_nent,
--        nent1=>AS_L1PHIHn1_AV_dout_nent,
--        nent2=>AS_L1PHIHn1_AV_dout_nent,
--        nent3=>AS_L1PHIHn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L1PHIHn1_V_readaddr
--      );

    AS_L1PHIHn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIHn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIHn1_wea_delay,
        addra     => AS_L1PHIHn1_writeaddr_delay,
        dina      => AS_L1PHIHn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIHn1_V_readaddr,
        doutb     => AS_L1PHIHn1_V_dout,
        sync_nent => AS_L1PHIHn1_start,
        nent_o    => AS_L1PHIHn1_AV_dout_nent
      );

    AS_L1PHIHn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIHn1_wea,
        addra     => AS_L1PHIHn1_writeaddr,
        dina      => AS_L1PHIHn1_din,
        wea_out       => AS_L1PHIHn1_wea_delay,
        addra_out     => AS_L1PHIHn1_writeaddr_delay,
        dina_out      => AS_L1PHIHn1_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIHn1_start
      );

    AS_L2PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L2PHIAn1_bx,
        bx_vld => AS_L2PHIAn1_bx_vld
      );

--    STREAM_AS_L2PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L2PHIAn1_bx,
--        bx_in_vld => AS_L2PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L2PHIAn1_stream_V_dout,
--        din0=>AS_L2PHIAn1_V_dout,
--        din1=>AS_L2PHIAn1_V_dout,
--        din2=>AS_L2PHIAn1_V_dout,
--        din3=>AS_L2PHIAn1_V_dout,
--        nent0=>AS_L2PHIAn1_AV_dout_nent,
--        nent1=>AS_L2PHIAn1_AV_dout_nent,
--        nent2=>AS_L2PHIAn1_AV_dout_nent,
--        nent3=>AS_L2PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L2PHIAn1_V_readaddr
--      );

    AS_L2PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIAn1_wea_delay,
        addra     => AS_L2PHIAn1_writeaddr_delay,
        dina      => AS_L2PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIAn1_V_readaddr,
        doutb     => AS_L2PHIAn1_V_dout,
        sync_nent => AS_L2PHIAn1_start,
        nent_o    => AS_L2PHIAn1_AV_dout_nent
      );

    AS_L2PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIAn1_wea,
        addra     => AS_L2PHIAn1_writeaddr,
        dina      => AS_L2PHIAn1_din,
        wea_out       => AS_L2PHIAn1_wea_delay,
        addra_out     => AS_L2PHIAn1_writeaddr_delay,
        dina_out      => AS_L2PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIAn1_start
      );

    AS_L2PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L2PHIBn1_bx,
        bx_vld => AS_L2PHIBn1_bx_vld
      );

--    STREAM_AS_L2PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L2PHIBn1_bx,
--        bx_in_vld => AS_L2PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L2PHIBn1_stream_V_dout,
--        din0=>AS_L2PHIBn1_V_dout,
--        din1=>AS_L2PHIBn1_V_dout,
--        din2=>AS_L2PHIBn1_V_dout,
--        din3=>AS_L2PHIBn1_V_dout,
--        nent0=>AS_L2PHIBn1_AV_dout_nent,
--        nent1=>AS_L2PHIBn1_AV_dout_nent,
--        nent2=>AS_L2PHIBn1_AV_dout_nent,
--        nent3=>AS_L2PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L2PHIBn1_V_readaddr
--      );

    AS_L2PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIBn1_wea_delay,
        addra     => AS_L2PHIBn1_writeaddr_delay,
        dina      => AS_L2PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIBn1_V_readaddr,
        doutb     => AS_L2PHIBn1_V_dout,
        sync_nent => AS_L2PHIBn1_start,
        nent_o    => AS_L2PHIBn1_AV_dout_nent
      );

    AS_L2PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIBn1_wea,
        addra     => AS_L2PHIBn1_writeaddr,
        dina      => AS_L2PHIBn1_din,
        wea_out       => AS_L2PHIBn1_wea_delay,
        addra_out     => AS_L2PHIBn1_writeaddr_delay,
        dina_out      => AS_L2PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIBn1_start
      );

    AS_L2PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L2PHICn1_bx,
        bx_vld => AS_L2PHICn1_bx_vld
      );

--    STREAM_AS_L2PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L2PHICn1_bx,
--        bx_in_vld => AS_L2PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L2PHICn1_stream_V_dout,
--        din0=>AS_L2PHICn1_V_dout,
--        din1=>AS_L2PHICn1_V_dout,
--        din2=>AS_L2PHICn1_V_dout,
--        din3=>AS_L2PHICn1_V_dout,
--        nent0=>AS_L2PHICn1_AV_dout_nent,
--        nent1=>AS_L2PHICn1_AV_dout_nent,
--        nent2=>AS_L2PHICn1_AV_dout_nent,
--        nent3=>AS_L2PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L2PHICn1_V_readaddr
--      );

    AS_L2PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHICn1_wea_delay,
        addra     => AS_L2PHICn1_writeaddr_delay,
        dina      => AS_L2PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHICn1_V_readaddr,
        doutb     => AS_L2PHICn1_V_dout,
        sync_nent => AS_L2PHICn1_start,
        nent_o    => AS_L2PHICn1_AV_dout_nent
      );

    AS_L2PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHICn1_wea,
        addra     => AS_L2PHICn1_writeaddr,
        dina      => AS_L2PHICn1_din,
        wea_out       => AS_L2PHICn1_wea_delay,
        addra_out     => AS_L2PHICn1_writeaddr_delay,
        dina_out      => AS_L2PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_L2PHICn1_start
      );

    AS_L2PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L2PHIDn1_bx,
        bx_vld => AS_L2PHIDn1_bx_vld
      );

--    STREAM_AS_L2PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L2PHIDn1_bx,
--        bx_in_vld => AS_L2PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L2PHIDn1_stream_V_dout,
--        din0=>AS_L2PHIDn1_V_dout,
--        din1=>AS_L2PHIDn1_V_dout,
--        din2=>AS_L2PHIDn1_V_dout,
--        din3=>AS_L2PHIDn1_V_dout,
--        nent0=>AS_L2PHIDn1_AV_dout_nent,
--        nent1=>AS_L2PHIDn1_AV_dout_nent,
--        nent2=>AS_L2PHIDn1_AV_dout_nent,
--        nent3=>AS_L2PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L2PHIDn1_V_readaddr
--      );

    AS_L2PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIDn1_wea_delay,
        addra     => AS_L2PHIDn1_writeaddr_delay,
        dina      => AS_L2PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIDn1_V_readaddr,
        doutb     => AS_L2PHIDn1_V_dout,
        sync_nent => AS_L2PHIDn1_start,
        nent_o    => AS_L2PHIDn1_AV_dout_nent
      );

    AS_L2PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIDn1_wea,
        addra     => AS_L2PHIDn1_writeaddr,
        dina      => AS_L2PHIDn1_din,
        wea_out       => AS_L2PHIDn1_wea_delay,
        addra_out     => AS_L2PHIDn1_writeaddr_delay,
        dina_out      => AS_L2PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIDn1_start
      );

    AS_L3PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L3PHIAn1_bx,
        bx_vld => AS_L3PHIAn1_bx_vld
      );

--    STREAM_AS_L3PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L3PHIAn1_bx,
--        bx_in_vld => AS_L3PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L3PHIAn1_stream_V_dout,
--        din0=>AS_L3PHIAn1_V_dout,
--        din1=>AS_L3PHIAn1_V_dout,
--        din2=>AS_L3PHIAn1_V_dout,
--        din3=>AS_L3PHIAn1_V_dout,
--        nent0=>AS_L3PHIAn1_AV_dout_nent,
--        nent1=>AS_L3PHIAn1_AV_dout_nent,
--        nent2=>AS_L3PHIAn1_AV_dout_nent,
--        nent3=>AS_L3PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L3PHIAn1_V_readaddr
--      );

    AS_L3PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIAn1_wea_delay,
        addra     => AS_L3PHIAn1_writeaddr_delay,
        dina      => AS_L3PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIAn1_V_readaddr,
        doutb     => AS_L3PHIAn1_V_dout,
        sync_nent => AS_L3PHIAn1_start,
        nent_o    => AS_L3PHIAn1_AV_dout_nent
      );

    AS_L3PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIAn1_wea,
        addra     => AS_L3PHIAn1_writeaddr,
        dina      => AS_L3PHIAn1_din,
        wea_out       => AS_L3PHIAn1_wea_delay,
        addra_out     => AS_L3PHIAn1_writeaddr_delay,
        dina_out      => AS_L3PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIAn1_start
      );

    AS_L3PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L3PHIBn1_bx,
        bx_vld => AS_L3PHIBn1_bx_vld
      );

--    STREAM_AS_L3PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L3PHIBn1_bx,
--        bx_in_vld => AS_L3PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L3PHIBn1_stream_V_dout,
--        din0=>AS_L3PHIBn1_V_dout,
--        din1=>AS_L3PHIBn1_V_dout,
--        din2=>AS_L3PHIBn1_V_dout,
--        din3=>AS_L3PHIBn1_V_dout,
--        nent0=>AS_L3PHIBn1_AV_dout_nent,
--        nent1=>AS_L3PHIBn1_AV_dout_nent,
--        nent2=>AS_L3PHIBn1_AV_dout_nent,
--        nent3=>AS_L3PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L3PHIBn1_V_readaddr
--      );

    AS_L3PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIBn1_wea_delay,
        addra     => AS_L3PHIBn1_writeaddr_delay,
        dina      => AS_L3PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIBn1_V_readaddr,
        doutb     => AS_L3PHIBn1_V_dout,
        sync_nent => AS_L3PHIBn1_start,
        nent_o    => AS_L3PHIBn1_AV_dout_nent
      );

    AS_L3PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIBn1_wea,
        addra     => AS_L3PHIBn1_writeaddr,
        dina      => AS_L3PHIBn1_din,
        wea_out       => AS_L3PHIBn1_wea_delay,
        addra_out     => AS_L3PHIBn1_writeaddr_delay,
        dina_out      => AS_L3PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIBn1_start
      );

    AS_L3PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L3PHICn1_bx,
        bx_vld => AS_L3PHICn1_bx_vld
      );

--    STREAM_AS_L3PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L3PHICn1_bx,
--        bx_in_vld => AS_L3PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L3PHICn1_stream_V_dout,
--        din0=>AS_L3PHICn1_V_dout,
--        din1=>AS_L3PHICn1_V_dout,
--        din2=>AS_L3PHICn1_V_dout,
--        din3=>AS_L3PHICn1_V_dout,
--        nent0=>AS_L3PHICn1_AV_dout_nent,
--        nent1=>AS_L3PHICn1_AV_dout_nent,
--        nent2=>AS_L3PHICn1_AV_dout_nent,
--        nent3=>AS_L3PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L3PHICn1_V_readaddr
--      );

    AS_L3PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHICn1_wea_delay,
        addra     => AS_L3PHICn1_writeaddr_delay,
        dina      => AS_L3PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHICn1_V_readaddr,
        doutb     => AS_L3PHICn1_V_dout,
        sync_nent => AS_L3PHICn1_start,
        nent_o    => AS_L3PHICn1_AV_dout_nent
      );

    AS_L3PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHICn1_wea,
        addra     => AS_L3PHICn1_writeaddr,
        dina      => AS_L3PHICn1_din,
        wea_out       => AS_L3PHICn1_wea_delay,
        addra_out     => AS_L3PHICn1_writeaddr_delay,
        dina_out      => AS_L3PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_L3PHICn1_start
      );

    AS_L3PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L3PHIDn1_bx,
        bx_vld => AS_L3PHIDn1_bx_vld
      );

--    STREAM_AS_L3PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L3PHIDn1_bx,
--        bx_in_vld => AS_L3PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L3PHIDn1_stream_V_dout,
--        din0=>AS_L3PHIDn1_V_dout,
--        din1=>AS_L3PHIDn1_V_dout,
--        din2=>AS_L3PHIDn1_V_dout,
--        din3=>AS_L3PHIDn1_V_dout,
--        nent0=>AS_L3PHIDn1_AV_dout_nent,
--        nent1=>AS_L3PHIDn1_AV_dout_nent,
--        nent2=>AS_L3PHIDn1_AV_dout_nent,
--        nent3=>AS_L3PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L3PHIDn1_V_readaddr
--      );

    AS_L3PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIDn1_wea_delay,
        addra     => AS_L3PHIDn1_writeaddr_delay,
        dina      => AS_L3PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIDn1_V_readaddr,
        doutb     => AS_L3PHIDn1_V_dout,
        sync_nent => AS_L3PHIDn1_start,
        nent_o    => AS_L3PHIDn1_AV_dout_nent
      );

    AS_L3PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIDn1_wea,
        addra     => AS_L3PHIDn1_writeaddr,
        dina      => AS_L3PHIDn1_din,
        wea_out       => AS_L3PHIDn1_wea_delay,
        addra_out     => AS_L3PHIDn1_writeaddr_delay,
        dina_out      => AS_L3PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIDn1_start
      );

    AS_L4PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L4PHIAn1_bx,
        bx_vld => AS_L4PHIAn1_bx_vld
      );

--    STREAM_AS_L4PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L4PHIAn1_bx,
--        bx_in_vld => AS_L4PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L4PHIAn1_stream_V_dout,
--        din0=>AS_L4PHIAn1_V_dout,
--        din1=>AS_L4PHIAn1_V_dout,
--        din2=>AS_L4PHIAn1_V_dout,
--        din3=>AS_L4PHIAn1_V_dout,
--        nent0=>AS_L4PHIAn1_AV_dout_nent,
--        nent1=>AS_L4PHIAn1_AV_dout_nent,
--        nent2=>AS_L4PHIAn1_AV_dout_nent,
--        nent3=>AS_L4PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L4PHIAn1_V_readaddr
--      );

    AS_L4PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIAn1_wea_delay,
        addra     => AS_L4PHIAn1_writeaddr_delay,
        dina      => AS_L4PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIAn1_V_readaddr,
        doutb     => AS_L4PHIAn1_V_dout,
        sync_nent => AS_L4PHIAn1_start,
        nent_o    => AS_L4PHIAn1_AV_dout_nent
      );

    AS_L4PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIAn1_wea,
        addra     => AS_L4PHIAn1_writeaddr,
        dina      => AS_L4PHIAn1_din,
        wea_out       => AS_L4PHIAn1_wea_delay,
        addra_out     => AS_L4PHIAn1_writeaddr_delay,
        dina_out      => AS_L4PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_L4PHIAn1_start
      );

    AS_L4PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L4PHIBn1_bx,
        bx_vld => AS_L4PHIBn1_bx_vld
      );

--    STREAM_AS_L4PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L4PHIBn1_bx,
--        bx_in_vld => AS_L4PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L4PHIBn1_stream_V_dout,
--        din0=>AS_L4PHIBn1_V_dout,
--        din1=>AS_L4PHIBn1_V_dout,
--        din2=>AS_L4PHIBn1_V_dout,
--        din3=>AS_L4PHIBn1_V_dout,
--        nent0=>AS_L4PHIBn1_AV_dout_nent,
--        nent1=>AS_L4PHIBn1_AV_dout_nent,
--        nent2=>AS_L4PHIBn1_AV_dout_nent,
--        nent3=>AS_L4PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L4PHIBn1_V_readaddr
--      );

    AS_L4PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIBn1_wea_delay,
        addra     => AS_L4PHIBn1_writeaddr_delay,
        dina      => AS_L4PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIBn1_V_readaddr,
        doutb     => AS_L4PHIBn1_V_dout,
        sync_nent => AS_L4PHIBn1_start,
        nent_o    => AS_L4PHIBn1_AV_dout_nent
      );

    AS_L4PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIBn1_wea,
        addra     => AS_L4PHIBn1_writeaddr,
        dina      => AS_L4PHIBn1_din,
        wea_out       => AS_L4PHIBn1_wea_delay,
        addra_out     => AS_L4PHIBn1_writeaddr_delay,
        dina_out      => AS_L4PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_L4PHIBn1_start
      );

    AS_L4PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L4PHICn1_bx,
        bx_vld => AS_L4PHICn1_bx_vld
      );

--    STREAM_AS_L4PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L4PHICn1_bx,
--        bx_in_vld => AS_L4PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L4PHICn1_stream_V_dout,
--        din0=>AS_L4PHICn1_V_dout,
--        din1=>AS_L4PHICn1_V_dout,
--        din2=>AS_L4PHICn1_V_dout,
--        din3=>AS_L4PHICn1_V_dout,
--        nent0=>AS_L4PHICn1_AV_dout_nent,
--        nent1=>AS_L4PHICn1_AV_dout_nent,
--        nent2=>AS_L4PHICn1_AV_dout_nent,
--        nent3=>AS_L4PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L4PHICn1_V_readaddr
--      );

    AS_L4PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHICn1_wea_delay,
        addra     => AS_L4PHICn1_writeaddr_delay,
        dina      => AS_L4PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHICn1_V_readaddr,
        doutb     => AS_L4PHICn1_V_dout,
        sync_nent => AS_L4PHICn1_start,
        nent_o    => AS_L4PHICn1_AV_dout_nent
      );

    AS_L4PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHICn1_wea,
        addra     => AS_L4PHICn1_writeaddr,
        dina      => AS_L4PHICn1_din,
        wea_out       => AS_L4PHICn1_wea_delay,
        addra_out     => AS_L4PHICn1_writeaddr_delay,
        dina_out      => AS_L4PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_L4PHICn1_start
      );

    AS_L4PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L4PHIDn1_bx,
        bx_vld => AS_L4PHIDn1_bx_vld
      );

--    STREAM_AS_L4PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L4PHIDn1_bx,
--        bx_in_vld => AS_L4PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L4PHIDn1_stream_V_dout,
--        din0=>AS_L4PHIDn1_V_dout,
--        din1=>AS_L4PHIDn1_V_dout,
--        din2=>AS_L4PHIDn1_V_dout,
--        din3=>AS_L4PHIDn1_V_dout,
--        nent0=>AS_L4PHIDn1_AV_dout_nent,
--        nent1=>AS_L4PHIDn1_AV_dout_nent,
--        nent2=>AS_L4PHIDn1_AV_dout_nent,
--        nent3=>AS_L4PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L4PHIDn1_V_readaddr
--      );

    AS_L4PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIDn1_wea_delay,
        addra     => AS_L4PHIDn1_writeaddr_delay,
        dina      => AS_L4PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIDn1_V_readaddr,
        doutb     => AS_L4PHIDn1_V_dout,
        sync_nent => AS_L4PHIDn1_start,
        nent_o    => AS_L4PHIDn1_AV_dout_nent
      );

    AS_L4PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIDn1_wea,
        addra     => AS_L4PHIDn1_writeaddr,
        dina      => AS_L4PHIDn1_din,
        wea_out       => AS_L4PHIDn1_wea_delay,
        addra_out     => AS_L4PHIDn1_writeaddr_delay,
        dina_out      => AS_L4PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_L4PHIDn1_start
      );

    AS_L5PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L5PHIAn1_bx,
        bx_vld => AS_L5PHIAn1_bx_vld
      );

--    STREAM_AS_L5PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L5PHIAn1_bx,
--        bx_in_vld => AS_L5PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L5PHIAn1_stream_V_dout,
--        din0=>AS_L5PHIAn1_V_dout,
--        din1=>AS_L5PHIAn1_V_dout,
--        din2=>AS_L5PHIAn1_V_dout,
--        din3=>AS_L5PHIAn1_V_dout,
--        nent0=>AS_L5PHIAn1_AV_dout_nent,
--        nent1=>AS_L5PHIAn1_AV_dout_nent,
--        nent2=>AS_L5PHIAn1_AV_dout_nent,
--        nent3=>AS_L5PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L5PHIAn1_V_readaddr
--      );

    AS_L5PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIAn1_wea_delay,
        addra     => AS_L5PHIAn1_writeaddr_delay,
        dina      => AS_L5PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIAn1_V_readaddr,
        doutb     => AS_L5PHIAn1_V_dout,
        sync_nent => AS_L5PHIAn1_start,
        nent_o    => AS_L5PHIAn1_AV_dout_nent
      );

    AS_L5PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIAn1_wea,
        addra     => AS_L5PHIAn1_writeaddr,
        dina      => AS_L5PHIAn1_din,
        wea_out       => AS_L5PHIAn1_wea_delay,
        addra_out     => AS_L5PHIAn1_writeaddr_delay,
        dina_out      => AS_L5PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIAn1_start
      );

    AS_L5PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L5PHIBn1_bx,
        bx_vld => AS_L5PHIBn1_bx_vld
      );

--    STREAM_AS_L5PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L5PHIBn1_bx,
--        bx_in_vld => AS_L5PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L5PHIBn1_stream_V_dout,
--        din0=>AS_L5PHIBn1_V_dout,
--        din1=>AS_L5PHIBn1_V_dout,
--        din2=>AS_L5PHIBn1_V_dout,
--        din3=>AS_L5PHIBn1_V_dout,
--        nent0=>AS_L5PHIBn1_AV_dout_nent,
--        nent1=>AS_L5PHIBn1_AV_dout_nent,
--        nent2=>AS_L5PHIBn1_AV_dout_nent,
--        nent3=>AS_L5PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L5PHIBn1_V_readaddr
--      );

    AS_L5PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIBn1_wea_delay,
        addra     => AS_L5PHIBn1_writeaddr_delay,
        dina      => AS_L5PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIBn1_V_readaddr,
        doutb     => AS_L5PHIBn1_V_dout,
        sync_nent => AS_L5PHIBn1_start,
        nent_o    => AS_L5PHIBn1_AV_dout_nent
      );

    AS_L5PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIBn1_wea,
        addra     => AS_L5PHIBn1_writeaddr,
        dina      => AS_L5PHIBn1_din,
        wea_out       => AS_L5PHIBn1_wea_delay,
        addra_out     => AS_L5PHIBn1_writeaddr_delay,
        dina_out      => AS_L5PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIBn1_start
      );

    AS_L5PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L5PHICn1_bx,
        bx_vld => AS_L5PHICn1_bx_vld
      );

--    STREAM_AS_L5PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L5PHICn1_bx,
--        bx_in_vld => AS_L5PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L5PHICn1_stream_V_dout,
--        din0=>AS_L5PHICn1_V_dout,
--        din1=>AS_L5PHICn1_V_dout,
--        din2=>AS_L5PHICn1_V_dout,
--        din3=>AS_L5PHICn1_V_dout,
--        nent0=>AS_L5PHICn1_AV_dout_nent,
--        nent1=>AS_L5PHICn1_AV_dout_nent,
--        nent2=>AS_L5PHICn1_AV_dout_nent,
--        nent3=>AS_L5PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L5PHICn1_V_readaddr
--      );

    AS_L5PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHICn1_wea_delay,
        addra     => AS_L5PHICn1_writeaddr_delay,
        dina      => AS_L5PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHICn1_V_readaddr,
        doutb     => AS_L5PHICn1_V_dout,
        sync_nent => AS_L5PHICn1_start,
        nent_o    => AS_L5PHICn1_AV_dout_nent
      );

    AS_L5PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHICn1_wea,
        addra     => AS_L5PHICn1_writeaddr,
        dina      => AS_L5PHICn1_din,
        wea_out       => AS_L5PHICn1_wea_delay,
        addra_out     => AS_L5PHICn1_writeaddr_delay,
        dina_out      => AS_L5PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_L5PHICn1_start
      );

    AS_L5PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L5PHIDn1_bx,
        bx_vld => AS_L5PHIDn1_bx_vld
      );

--    STREAM_AS_L5PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L5PHIDn1_bx,
--        bx_in_vld => AS_L5PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L5PHIDn1_stream_V_dout,
--        din0=>AS_L5PHIDn1_V_dout,
--        din1=>AS_L5PHIDn1_V_dout,
--        din2=>AS_L5PHIDn1_V_dout,
--        din3=>AS_L5PHIDn1_V_dout,
--        nent0=>AS_L5PHIDn1_AV_dout_nent,
--        nent1=>AS_L5PHIDn1_AV_dout_nent,
--        nent2=>AS_L5PHIDn1_AV_dout_nent,
--        nent3=>AS_L5PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L5PHIDn1_V_readaddr
--      );

    AS_L5PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIDn1_wea_delay,
        addra     => AS_L5PHIDn1_writeaddr_delay,
        dina      => AS_L5PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIDn1_V_readaddr,
        doutb     => AS_L5PHIDn1_V_dout,
        sync_nent => AS_L5PHIDn1_start,
        nent_o    => AS_L5PHIDn1_AV_dout_nent
      );

    AS_L5PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIDn1_wea,
        addra     => AS_L5PHIDn1_writeaddr,
        dina      => AS_L5PHIDn1_din,
        wea_out       => AS_L5PHIDn1_wea_delay,
        addra_out     => AS_L5PHIDn1_writeaddr_delay,
        dina_out      => AS_L5PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIDn1_start
      );

    AS_L6PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L6PHIAn1_bx,
        bx_vld => AS_L6PHIAn1_bx_vld
      );

--    STREAM_AS_L6PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L6PHIAn1_bx,
--        bx_in_vld => AS_L6PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L6PHIAn1_stream_V_dout,
--        din0=>AS_L6PHIAn1_V_dout,
--        din1=>AS_L6PHIAn1_V_dout,
--        din2=>AS_L6PHIAn1_V_dout,
--        din3=>AS_L6PHIAn1_V_dout,
--        nent0=>AS_L6PHIAn1_AV_dout_nent,
--        nent1=>AS_L6PHIAn1_AV_dout_nent,
--        nent2=>AS_L6PHIAn1_AV_dout_nent,
--        nent3=>AS_L6PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L6PHIAn1_V_readaddr
--      );

    AS_L6PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIAn1_wea_delay,
        addra     => AS_L6PHIAn1_writeaddr_delay,
        dina      => AS_L6PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIAn1_V_readaddr,
        doutb     => AS_L6PHIAn1_V_dout,
        sync_nent => AS_L6PHIAn1_start,
        nent_o    => AS_L6PHIAn1_AV_dout_nent
      );

    AS_L6PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIAn1_wea,
        addra     => AS_L6PHIAn1_writeaddr,
        dina      => AS_L6PHIAn1_din,
        wea_out       => AS_L6PHIAn1_wea_delay,
        addra_out     => AS_L6PHIAn1_writeaddr_delay,
        dina_out      => AS_L6PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_L6PHIAn1_start
      );

    AS_L6PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L6PHIBn1_bx,
        bx_vld => AS_L6PHIBn1_bx_vld
      );

--    STREAM_AS_L6PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L6PHIBn1_bx,
--        bx_in_vld => AS_L6PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L6PHIBn1_stream_V_dout,
--        din0=>AS_L6PHIBn1_V_dout,
--        din1=>AS_L6PHIBn1_V_dout,
--        din2=>AS_L6PHIBn1_V_dout,
--        din3=>AS_L6PHIBn1_V_dout,
--        nent0=>AS_L6PHIBn1_AV_dout_nent,
--        nent1=>AS_L6PHIBn1_AV_dout_nent,
--        nent2=>AS_L6PHIBn1_AV_dout_nent,
--        nent3=>AS_L6PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L6PHIBn1_V_readaddr
--      );

    AS_L6PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIBn1_wea_delay,
        addra     => AS_L6PHIBn1_writeaddr_delay,
        dina      => AS_L6PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIBn1_V_readaddr,
        doutb     => AS_L6PHIBn1_V_dout,
        sync_nent => AS_L6PHIBn1_start,
        nent_o    => AS_L6PHIBn1_AV_dout_nent
      );

    AS_L6PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIBn1_wea,
        addra     => AS_L6PHIBn1_writeaddr,
        dina      => AS_L6PHIBn1_din,
        wea_out       => AS_L6PHIBn1_wea_delay,
        addra_out     => AS_L6PHIBn1_writeaddr_delay,
        dina_out      => AS_L6PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_L6PHIBn1_start
      );

    AS_L6PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L6PHICn1_bx,
        bx_vld => AS_L6PHICn1_bx_vld
      );

--    STREAM_AS_L6PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L6PHICn1_bx,
--        bx_in_vld => AS_L6PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L6PHICn1_stream_V_dout,
--        din0=>AS_L6PHICn1_V_dout,
--        din1=>AS_L6PHICn1_V_dout,
--        din2=>AS_L6PHICn1_V_dout,
--        din3=>AS_L6PHICn1_V_dout,
--        nent0=>AS_L6PHICn1_AV_dout_nent,
--        nent1=>AS_L6PHICn1_AV_dout_nent,
--        nent2=>AS_L6PHICn1_AV_dout_nent,
--        nent3=>AS_L6PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L6PHICn1_V_readaddr
--      );

    AS_L6PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHICn1_wea_delay,
        addra     => AS_L6PHICn1_writeaddr_delay,
        dina      => AS_L6PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHICn1_V_readaddr,
        doutb     => AS_L6PHICn1_V_dout,
        sync_nent => AS_L6PHICn1_start,
        nent_o    => AS_L6PHICn1_AV_dout_nent
      );

    AS_L6PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHICn1_wea,
        addra     => AS_L6PHICn1_writeaddr,
        dina      => AS_L6PHICn1_din,
        wea_out       => AS_L6PHICn1_wea_delay,
        addra_out     => AS_L6PHICn1_writeaddr_delay,
        dina_out      => AS_L6PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_L6PHICn1_start
      );

    AS_L6PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_L6PHIDn1_bx,
        bx_vld => AS_L6PHIDn1_bx_vld
      );

--    STREAM_AS_L6PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_L6PHIDn1_bx,
--        bx_in_vld => AS_L6PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_L6PHIDn1_stream_V_dout,
--        din0=>AS_L6PHIDn1_V_dout,
--        din1=>AS_L6PHIDn1_V_dout,
--        din2=>AS_L6PHIDn1_V_dout,
--        din3=>AS_L6PHIDn1_V_dout,
--        nent0=>AS_L6PHIDn1_AV_dout_nent,
--        nent1=>AS_L6PHIDn1_AV_dout_nent,
--        nent2=>AS_L6PHIDn1_AV_dout_nent,
--        nent3=>AS_L6PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_L6PHIDn1_V_readaddr
--      );

    AS_L6PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIDn1_wea_delay,
        addra     => AS_L6PHIDn1_writeaddr_delay,
        dina      => AS_L6PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIDn1_V_readaddr,
        doutb     => AS_L6PHIDn1_V_dout,
        sync_nent => AS_L6PHIDn1_start,
        nent_o    => AS_L6PHIDn1_AV_dout_nent
      );

    AS_L6PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIDn1_wea,
        addra     => AS_L6PHIDn1_writeaddr,
        dina      => AS_L6PHIDn1_din,
        wea_out       => AS_L6PHIDn1_wea_delay,
        addra_out     => AS_L6PHIDn1_writeaddr_delay,
        dina_out      => AS_L6PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_L6PHIDn1_start
      );

    AS_D1PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D1PHIAn1_bx,
        bx_vld => AS_D1PHIAn1_bx_vld
      );

--    STREAM_AS_D1PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D1PHIAn1_bx,
--        bx_in_vld => AS_D1PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D1PHIAn1_stream_V_dout,
--        din0=>AS_D1PHIAn1_V_dout,
--        din1=>AS_D1PHIAn1_V_dout,
--        din2=>AS_D1PHIAn1_V_dout,
--        din3=>AS_D1PHIAn1_V_dout,
--        nent0=>AS_D1PHIAn1_AV_dout_nent,
--        nent1=>AS_D1PHIAn1_AV_dout_nent,
--        nent2=>AS_D1PHIAn1_AV_dout_nent,
--        nent3=>AS_D1PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D1PHIAn1_V_readaddr
--      );

    AS_D1PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIAn1_wea_delay,
        addra     => AS_D1PHIAn1_writeaddr_delay,
        dina      => AS_D1PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIAn1_V_readaddr,
        doutb     => AS_D1PHIAn1_V_dout,
        sync_nent => AS_D1PHIAn1_start,
        nent_o    => AS_D1PHIAn1_AV_dout_nent
      );

    AS_D1PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIAn1_wea,
        addra     => AS_D1PHIAn1_writeaddr,
        dina      => AS_D1PHIAn1_din,
        wea_out       => AS_D1PHIAn1_wea_delay,
        addra_out     => AS_D1PHIAn1_writeaddr_delay,
        dina_out      => AS_D1PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIAn1_start
      );

    AS_D1PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D1PHIBn1_bx,
        bx_vld => AS_D1PHIBn1_bx_vld
      );

--    STREAM_AS_D1PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D1PHIBn1_bx,
--        bx_in_vld => AS_D1PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D1PHIBn1_stream_V_dout,
--        din0=>AS_D1PHIBn1_V_dout,
--        din1=>AS_D1PHIBn1_V_dout,
--        din2=>AS_D1PHIBn1_V_dout,
--        din3=>AS_D1PHIBn1_V_dout,
--        nent0=>AS_D1PHIBn1_AV_dout_nent,
--        nent1=>AS_D1PHIBn1_AV_dout_nent,
--        nent2=>AS_D1PHIBn1_AV_dout_nent,
--        nent3=>AS_D1PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D1PHIBn1_V_readaddr
--      );

    AS_D1PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIBn1_wea_delay,
        addra     => AS_D1PHIBn1_writeaddr_delay,
        dina      => AS_D1PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIBn1_V_readaddr,
        doutb     => AS_D1PHIBn1_V_dout,
        sync_nent => AS_D1PHIBn1_start,
        nent_o    => AS_D1PHIBn1_AV_dout_nent
      );

    AS_D1PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIBn1_wea,
        addra     => AS_D1PHIBn1_writeaddr,
        dina      => AS_D1PHIBn1_din,
        wea_out       => AS_D1PHIBn1_wea_delay,
        addra_out     => AS_D1PHIBn1_writeaddr_delay,
        dina_out      => AS_D1PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIBn1_start
      );

    AS_D1PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D1PHICn1_bx,
        bx_vld => AS_D1PHICn1_bx_vld
      );

--    STREAM_AS_D1PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D1PHICn1_bx,
--        bx_in_vld => AS_D1PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D1PHICn1_stream_V_dout,
--        din0=>AS_D1PHICn1_V_dout,
--        din1=>AS_D1PHICn1_V_dout,
--        din2=>AS_D1PHICn1_V_dout,
--        din3=>AS_D1PHICn1_V_dout,
--        nent0=>AS_D1PHICn1_AV_dout_nent,
--        nent1=>AS_D1PHICn1_AV_dout_nent,
--        nent2=>AS_D1PHICn1_AV_dout_nent,
--        nent3=>AS_D1PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D1PHICn1_V_readaddr
--      );

    AS_D1PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHICn1_wea_delay,
        addra     => AS_D1PHICn1_writeaddr_delay,
        dina      => AS_D1PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHICn1_V_readaddr,
        doutb     => AS_D1PHICn1_V_dout,
        sync_nent => AS_D1PHICn1_start,
        nent_o    => AS_D1PHICn1_AV_dout_nent
      );

    AS_D1PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHICn1_wea,
        addra     => AS_D1PHICn1_writeaddr,
        dina      => AS_D1PHICn1_din,
        wea_out       => AS_D1PHICn1_wea_delay,
        addra_out     => AS_D1PHICn1_writeaddr_delay,
        dina_out      => AS_D1PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_D1PHICn1_start
      );

    AS_D1PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D1PHIDn1_bx,
        bx_vld => AS_D1PHIDn1_bx_vld
      );

--    STREAM_AS_D1PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D1PHIDn1_bx,
--        bx_in_vld => AS_D1PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D1PHIDn1_stream_V_dout,
--        din0=>AS_D1PHIDn1_V_dout,
--        din1=>AS_D1PHIDn1_V_dout,
--        din2=>AS_D1PHIDn1_V_dout,
--        din3=>AS_D1PHIDn1_V_dout,
--        nent0=>AS_D1PHIDn1_AV_dout_nent,
--        nent1=>AS_D1PHIDn1_AV_dout_nent,
--        nent2=>AS_D1PHIDn1_AV_dout_nent,
--        nent3=>AS_D1PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D1PHIDn1_V_readaddr
--      );

    AS_D1PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIDn1_wea_delay,
        addra     => AS_D1PHIDn1_writeaddr_delay,
        dina      => AS_D1PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIDn1_V_readaddr,
        doutb     => AS_D1PHIDn1_V_dout,
        sync_nent => AS_D1PHIDn1_start,
        nent_o    => AS_D1PHIDn1_AV_dout_nent
      );

    AS_D1PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIDn1_wea,
        addra     => AS_D1PHIDn1_writeaddr,
        dina      => AS_D1PHIDn1_din,
        wea_out       => AS_D1PHIDn1_wea_delay,
        addra_out     => AS_D1PHIDn1_writeaddr_delay,
        dina_out      => AS_D1PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIDn1_start
      );

    AS_D2PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D2PHIAn1_bx,
        bx_vld => AS_D2PHIAn1_bx_vld
      );

--    STREAM_AS_D2PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D2PHIAn1_bx,
--        bx_in_vld => AS_D2PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D2PHIAn1_stream_V_dout,
--        din0=>AS_D2PHIAn1_V_dout,
--        din1=>AS_D2PHIAn1_V_dout,
--        din2=>AS_D2PHIAn1_V_dout,
--        din3=>AS_D2PHIAn1_V_dout,
--        nent0=>AS_D2PHIAn1_AV_dout_nent,
--        nent1=>AS_D2PHIAn1_AV_dout_nent,
--        nent2=>AS_D2PHIAn1_AV_dout_nent,
--        nent3=>AS_D2PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D2PHIAn1_V_readaddr
--      );

    AS_D2PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIAn1_wea_delay,
        addra     => AS_D2PHIAn1_writeaddr_delay,
        dina      => AS_D2PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIAn1_V_readaddr,
        doutb     => AS_D2PHIAn1_V_dout,
        sync_nent => AS_D2PHIAn1_start,
        nent_o    => AS_D2PHIAn1_AV_dout_nent
      );

    AS_D2PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIAn1_wea,
        addra     => AS_D2PHIAn1_writeaddr,
        dina      => AS_D2PHIAn1_din,
        wea_out       => AS_D2PHIAn1_wea_delay,
        addra_out     => AS_D2PHIAn1_writeaddr_delay,
        dina_out      => AS_D2PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_D2PHIAn1_start
      );

    AS_D2PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D2PHIBn1_bx,
        bx_vld => AS_D2PHIBn1_bx_vld
      );

--    STREAM_AS_D2PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D2PHIBn1_bx,
--        bx_in_vld => AS_D2PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D2PHIBn1_stream_V_dout,
--        din0=>AS_D2PHIBn1_V_dout,
--        din1=>AS_D2PHIBn1_V_dout,
--        din2=>AS_D2PHIBn1_V_dout,
--        din3=>AS_D2PHIBn1_V_dout,
--        nent0=>AS_D2PHIBn1_AV_dout_nent,
--        nent1=>AS_D2PHIBn1_AV_dout_nent,
--        nent2=>AS_D2PHIBn1_AV_dout_nent,
--        nent3=>AS_D2PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D2PHIBn1_V_readaddr
--      );

    AS_D2PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIBn1_wea_delay,
        addra     => AS_D2PHIBn1_writeaddr_delay,
        dina      => AS_D2PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIBn1_V_readaddr,
        doutb     => AS_D2PHIBn1_V_dout,
        sync_nent => AS_D2PHIBn1_start,
        nent_o    => AS_D2PHIBn1_AV_dout_nent
      );

    AS_D2PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIBn1_wea,
        addra     => AS_D2PHIBn1_writeaddr,
        dina      => AS_D2PHIBn1_din,
        wea_out       => AS_D2PHIBn1_wea_delay,
        addra_out     => AS_D2PHIBn1_writeaddr_delay,
        dina_out      => AS_D2PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_D2PHIBn1_start
      );

    AS_D2PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D2PHICn1_bx,
        bx_vld => AS_D2PHICn1_bx_vld
      );

--    STREAM_AS_D2PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D2PHICn1_bx,
--        bx_in_vld => AS_D2PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D2PHICn1_stream_V_dout,
--        din0=>AS_D2PHICn1_V_dout,
--        din1=>AS_D2PHICn1_V_dout,
--        din2=>AS_D2PHICn1_V_dout,
--        din3=>AS_D2PHICn1_V_dout,
--        nent0=>AS_D2PHICn1_AV_dout_nent,
--        nent1=>AS_D2PHICn1_AV_dout_nent,
--        nent2=>AS_D2PHICn1_AV_dout_nent,
--        nent3=>AS_D2PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D2PHICn1_V_readaddr
--      );

    AS_D2PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHICn1_wea_delay,
        addra     => AS_D2PHICn1_writeaddr_delay,
        dina      => AS_D2PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHICn1_V_readaddr,
        doutb     => AS_D2PHICn1_V_dout,
        sync_nent => AS_D2PHICn1_start,
        nent_o    => AS_D2PHICn1_AV_dout_nent
      );

    AS_D2PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHICn1_wea,
        addra     => AS_D2PHICn1_writeaddr,
        dina      => AS_D2PHICn1_din,
        wea_out       => AS_D2PHICn1_wea_delay,
        addra_out     => AS_D2PHICn1_writeaddr_delay,
        dina_out      => AS_D2PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_D2PHICn1_start
      );

    AS_D2PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D2PHIDn1_bx,
        bx_vld => AS_D2PHIDn1_bx_vld
      );

--    STREAM_AS_D2PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D2PHIDn1_bx,
--        bx_in_vld => AS_D2PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D2PHIDn1_stream_V_dout,
--        din0=>AS_D2PHIDn1_V_dout,
--        din1=>AS_D2PHIDn1_V_dout,
--        din2=>AS_D2PHIDn1_V_dout,
--        din3=>AS_D2PHIDn1_V_dout,
--        nent0=>AS_D2PHIDn1_AV_dout_nent,
--        nent1=>AS_D2PHIDn1_AV_dout_nent,
--        nent2=>AS_D2PHIDn1_AV_dout_nent,
--        nent3=>AS_D2PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D2PHIDn1_V_readaddr
--      );

    AS_D2PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIDn1_wea_delay,
        addra     => AS_D2PHIDn1_writeaddr_delay,
        dina      => AS_D2PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIDn1_V_readaddr,
        doutb     => AS_D2PHIDn1_V_dout,
        sync_nent => AS_D2PHIDn1_start,
        nent_o    => AS_D2PHIDn1_AV_dout_nent
      );

    AS_D2PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIDn1_wea,
        addra     => AS_D2PHIDn1_writeaddr,
        dina      => AS_D2PHIDn1_din,
        wea_out       => AS_D2PHIDn1_wea_delay,
        addra_out     => AS_D2PHIDn1_writeaddr_delay,
        dina_out      => AS_D2PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_D2PHIDn1_start
      );

    AS_D3PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D3PHIAn1_bx,
        bx_vld => AS_D3PHIAn1_bx_vld
      );

--    STREAM_AS_D3PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D3PHIAn1_bx,
--        bx_in_vld => AS_D3PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D3PHIAn1_stream_V_dout,
--        din0=>AS_D3PHIAn1_V_dout,
--        din1=>AS_D3PHIAn1_V_dout,
--        din2=>AS_D3PHIAn1_V_dout,
--        din3=>AS_D3PHIAn1_V_dout,
--        nent0=>AS_D3PHIAn1_AV_dout_nent,
--        nent1=>AS_D3PHIAn1_AV_dout_nent,
--        nent2=>AS_D3PHIAn1_AV_dout_nent,
--        nent3=>AS_D3PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D3PHIAn1_V_readaddr
--      );

    AS_D3PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIAn1_wea_delay,
        addra     => AS_D3PHIAn1_writeaddr_delay,
        dina      => AS_D3PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIAn1_V_readaddr,
        doutb     => AS_D3PHIAn1_V_dout,
        sync_nent => AS_D3PHIAn1_start,
        nent_o    => AS_D3PHIAn1_AV_dout_nent
      );

    AS_D3PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIAn1_wea,
        addra     => AS_D3PHIAn1_writeaddr,
        dina      => AS_D3PHIAn1_din,
        wea_out       => AS_D3PHIAn1_wea_delay,
        addra_out     => AS_D3PHIAn1_writeaddr_delay,
        dina_out      => AS_D3PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIAn1_start
      );

    AS_D3PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D3PHIBn1_bx,
        bx_vld => AS_D3PHIBn1_bx_vld
      );

--    STREAM_AS_D3PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D3PHIBn1_bx,
--        bx_in_vld => AS_D3PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D3PHIBn1_stream_V_dout,
--        din0=>AS_D3PHIBn1_V_dout,
--        din1=>AS_D3PHIBn1_V_dout,
--        din2=>AS_D3PHIBn1_V_dout,
--        din3=>AS_D3PHIBn1_V_dout,
--        nent0=>AS_D3PHIBn1_AV_dout_nent,
--        nent1=>AS_D3PHIBn1_AV_dout_nent,
--        nent2=>AS_D3PHIBn1_AV_dout_nent,
--        nent3=>AS_D3PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D3PHIBn1_V_readaddr
--      );

    AS_D3PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIBn1_wea_delay,
        addra     => AS_D3PHIBn1_writeaddr_delay,
        dina      => AS_D3PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIBn1_V_readaddr,
        doutb     => AS_D3PHIBn1_V_dout,
        sync_nent => AS_D3PHIBn1_start,
        nent_o    => AS_D3PHIBn1_AV_dout_nent
      );

    AS_D3PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIBn1_wea,
        addra     => AS_D3PHIBn1_writeaddr,
        dina      => AS_D3PHIBn1_din,
        wea_out       => AS_D3PHIBn1_wea_delay,
        addra_out     => AS_D3PHIBn1_writeaddr_delay,
        dina_out      => AS_D3PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIBn1_start
      );

    AS_D3PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D3PHICn1_bx,
        bx_vld => AS_D3PHICn1_bx_vld
      );

--    STREAM_AS_D3PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D3PHICn1_bx,
--        bx_in_vld => AS_D3PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D3PHICn1_stream_V_dout,
--        din0=>AS_D3PHICn1_V_dout,
--        din1=>AS_D3PHICn1_V_dout,
--        din2=>AS_D3PHICn1_V_dout,
--        din3=>AS_D3PHICn1_V_dout,
--        nent0=>AS_D3PHICn1_AV_dout_nent,
--        nent1=>AS_D3PHICn1_AV_dout_nent,
--        nent2=>AS_D3PHICn1_AV_dout_nent,
--        nent3=>AS_D3PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D3PHICn1_V_readaddr
--      );

    AS_D3PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHICn1_wea_delay,
        addra     => AS_D3PHICn1_writeaddr_delay,
        dina      => AS_D3PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHICn1_V_readaddr,
        doutb     => AS_D3PHICn1_V_dout,
        sync_nent => AS_D3PHICn1_start,
        nent_o    => AS_D3PHICn1_AV_dout_nent
      );

    AS_D3PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHICn1_wea,
        addra     => AS_D3PHICn1_writeaddr,
        dina      => AS_D3PHICn1_din,
        wea_out       => AS_D3PHICn1_wea_delay,
        addra_out     => AS_D3PHICn1_writeaddr_delay,
        dina_out      => AS_D3PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_D3PHICn1_start
      );

    AS_D3PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D3PHIDn1_bx,
        bx_vld => AS_D3PHIDn1_bx_vld
      );

--    STREAM_AS_D3PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D3PHIDn1_bx,
--        bx_in_vld => AS_D3PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D3PHIDn1_stream_V_dout,
--        din0=>AS_D3PHIDn1_V_dout,
--        din1=>AS_D3PHIDn1_V_dout,
--        din2=>AS_D3PHIDn1_V_dout,
--        din3=>AS_D3PHIDn1_V_dout,
--        nent0=>AS_D3PHIDn1_AV_dout_nent,
--        nent1=>AS_D3PHIDn1_AV_dout_nent,
--        nent2=>AS_D3PHIDn1_AV_dout_nent,
--        nent3=>AS_D3PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D3PHIDn1_V_readaddr
--      );

    AS_D3PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIDn1_wea_delay,
        addra     => AS_D3PHIDn1_writeaddr_delay,
        dina      => AS_D3PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIDn1_V_readaddr,
        doutb     => AS_D3PHIDn1_V_dout,
        sync_nent => AS_D3PHIDn1_start,
        nent_o    => AS_D3PHIDn1_AV_dout_nent
      );

    AS_D3PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIDn1_wea,
        addra     => AS_D3PHIDn1_writeaddr,
        dina      => AS_D3PHIDn1_din,
        wea_out       => AS_D3PHIDn1_wea_delay,
        addra_out     => AS_D3PHIDn1_writeaddr_delay,
        dina_out      => AS_D3PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIDn1_start
      );

    AS_D4PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D4PHIAn1_bx,
        bx_vld => AS_D4PHIAn1_bx_vld
      );

--    STREAM_AS_D4PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D4PHIAn1_bx,
--        bx_in_vld => AS_D4PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D4PHIAn1_stream_V_dout,
--        din0=>AS_D4PHIAn1_V_dout,
--        din1=>AS_D4PHIAn1_V_dout,
--        din2=>AS_D4PHIAn1_V_dout,
--        din3=>AS_D4PHIAn1_V_dout,
--        nent0=>AS_D4PHIAn1_AV_dout_nent,
--        nent1=>AS_D4PHIAn1_AV_dout_nent,
--        nent2=>AS_D4PHIAn1_AV_dout_nent,
--        nent3=>AS_D4PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D4PHIAn1_V_readaddr
--      );

    AS_D4PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIAn1_wea_delay,
        addra     => AS_D4PHIAn1_writeaddr_delay,
        dina      => AS_D4PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIAn1_V_readaddr,
        doutb     => AS_D4PHIAn1_V_dout,
        sync_nent => AS_D4PHIAn1_start,
        nent_o    => AS_D4PHIAn1_AV_dout_nent
      );

    AS_D4PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIAn1_wea,
        addra     => AS_D4PHIAn1_writeaddr,
        dina      => AS_D4PHIAn1_din,
        wea_out       => AS_D4PHIAn1_wea_delay,
        addra_out     => AS_D4PHIAn1_writeaddr_delay,
        dina_out      => AS_D4PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_D4PHIAn1_start
      );

    AS_D4PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D4PHIBn1_bx,
        bx_vld => AS_D4PHIBn1_bx_vld
      );

--    STREAM_AS_D4PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D4PHIBn1_bx,
--        bx_in_vld => AS_D4PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D4PHIBn1_stream_V_dout,
--        din0=>AS_D4PHIBn1_V_dout,
--        din1=>AS_D4PHIBn1_V_dout,
--        din2=>AS_D4PHIBn1_V_dout,
--        din3=>AS_D4PHIBn1_V_dout,
--        nent0=>AS_D4PHIBn1_AV_dout_nent,
--        nent1=>AS_D4PHIBn1_AV_dout_nent,
--        nent2=>AS_D4PHIBn1_AV_dout_nent,
--        nent3=>AS_D4PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D4PHIBn1_V_readaddr
--      );

    AS_D4PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIBn1_wea_delay,
        addra     => AS_D4PHIBn1_writeaddr_delay,
        dina      => AS_D4PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIBn1_V_readaddr,
        doutb     => AS_D4PHIBn1_V_dout,
        sync_nent => AS_D4PHIBn1_start,
        nent_o    => AS_D4PHIBn1_AV_dout_nent
      );

    AS_D4PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIBn1_wea,
        addra     => AS_D4PHIBn1_writeaddr,
        dina      => AS_D4PHIBn1_din,
        wea_out       => AS_D4PHIBn1_wea_delay,
        addra_out     => AS_D4PHIBn1_writeaddr_delay,
        dina_out      => AS_D4PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_D4PHIBn1_start
      );

    AS_D4PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D4PHICn1_bx,
        bx_vld => AS_D4PHICn1_bx_vld
      );

--    STREAM_AS_D4PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D4PHICn1_bx,
--        bx_in_vld => AS_D4PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D4PHICn1_stream_V_dout,
--        din0=>AS_D4PHICn1_V_dout,
--        din1=>AS_D4PHICn1_V_dout,
--        din2=>AS_D4PHICn1_V_dout,
--        din3=>AS_D4PHICn1_V_dout,
--        nent0=>AS_D4PHICn1_AV_dout_nent,
--        nent1=>AS_D4PHICn1_AV_dout_nent,
--        nent2=>AS_D4PHICn1_AV_dout_nent,
--        nent3=>AS_D4PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D4PHICn1_V_readaddr
--      );

    AS_D4PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHICn1_wea_delay,
        addra     => AS_D4PHICn1_writeaddr_delay,
        dina      => AS_D4PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHICn1_V_readaddr,
        doutb     => AS_D4PHICn1_V_dout,
        sync_nent => AS_D4PHICn1_start,
        nent_o    => AS_D4PHICn1_AV_dout_nent
      );

    AS_D4PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHICn1_wea,
        addra     => AS_D4PHICn1_writeaddr,
        dina      => AS_D4PHICn1_din,
        wea_out       => AS_D4PHICn1_wea_delay,
        addra_out     => AS_D4PHICn1_writeaddr_delay,
        dina_out      => AS_D4PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_D4PHICn1_start
      );

    AS_D4PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D4PHIDn1_bx,
        bx_vld => AS_D4PHIDn1_bx_vld
      );

--    STREAM_AS_D4PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D4PHIDn1_bx,
--        bx_in_vld => AS_D4PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D4PHIDn1_stream_V_dout,
--        din0=>AS_D4PHIDn1_V_dout,
--        din1=>AS_D4PHIDn1_V_dout,
--        din2=>AS_D4PHIDn1_V_dout,
--        din3=>AS_D4PHIDn1_V_dout,
--        nent0=>AS_D4PHIDn1_AV_dout_nent,
--        nent1=>AS_D4PHIDn1_AV_dout_nent,
--        nent2=>AS_D4PHIDn1_AV_dout_nent,
--        nent3=>AS_D4PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D4PHIDn1_V_readaddr
--      );

    AS_D4PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIDn1_wea_delay,
        addra     => AS_D4PHIDn1_writeaddr_delay,
        dina      => AS_D4PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIDn1_V_readaddr,
        doutb     => AS_D4PHIDn1_V_dout,
        sync_nent => AS_D4PHIDn1_start,
        nent_o    => AS_D4PHIDn1_AV_dout_nent
      );

    AS_D4PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIDn1_wea,
        addra     => AS_D4PHIDn1_writeaddr,
        dina      => AS_D4PHIDn1_din,
        wea_out       => AS_D4PHIDn1_wea_delay,
        addra_out     => AS_D4PHIDn1_writeaddr_delay,
        dina_out      => AS_D4PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_D4PHIDn1_start
      );

    AS_D5PHIAn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D5PHIAn1_bx,
        bx_vld => AS_D5PHIAn1_bx_vld
      );

--    STREAM_AS_D5PHIAn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D5PHIAn1_bx,
--        bx_in_vld => AS_D5PHIAn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D5PHIAn1_stream_V_dout,
--        din0=>AS_D5PHIAn1_V_dout,
--        din1=>AS_D5PHIAn1_V_dout,
--        din2=>AS_D5PHIAn1_V_dout,
--        din3=>AS_D5PHIAn1_V_dout,
--        nent0=>AS_D5PHIAn1_AV_dout_nent,
--        nent1=>AS_D5PHIAn1_AV_dout_nent,
--        nent2=>AS_D5PHIAn1_AV_dout_nent,
--        nent3=>AS_D5PHIAn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D5PHIAn1_V_readaddr
--      );

    AS_D5PHIAn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIAn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIAn1_wea_delay,
        addra     => AS_D5PHIAn1_writeaddr_delay,
        dina      => AS_D5PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIAn1_V_readaddr,
        doutb     => AS_D5PHIAn1_V_dout,
        sync_nent => AS_D5PHIAn1_start,
        nent_o    => AS_D5PHIAn1_AV_dout_nent
      );

    AS_D5PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIAn1_wea,
        addra     => AS_D5PHIAn1_writeaddr,
        dina      => AS_D5PHIAn1_din,
        wea_out       => AS_D5PHIAn1_wea_delay,
        addra_out     => AS_D5PHIAn1_writeaddr_delay,
        dina_out      => AS_D5PHIAn1_din_delay,
        done       => VMR_done,
        start      => AS_D5PHIAn1_start
      );

    AS_D5PHIBn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D5PHIBn1_bx,
        bx_vld => AS_D5PHIBn1_bx_vld
      );

--    STREAM_AS_D5PHIBn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D5PHIBn1_bx,
--        bx_in_vld => AS_D5PHIBn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D5PHIBn1_stream_V_dout,
--        din0=>AS_D5PHIBn1_V_dout,
--        din1=>AS_D5PHIBn1_V_dout,
--        din2=>AS_D5PHIBn1_V_dout,
--        din3=>AS_D5PHIBn1_V_dout,
--        nent0=>AS_D5PHIBn1_AV_dout_nent,
--        nent1=>AS_D5PHIBn1_AV_dout_nent,
--        nent2=>AS_D5PHIBn1_AV_dout_nent,
--        nent3=>AS_D5PHIBn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D5PHIBn1_V_readaddr
--      );

    AS_D5PHIBn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIBn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIBn1_wea_delay,
        addra     => AS_D5PHIBn1_writeaddr_delay,
        dina      => AS_D5PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIBn1_V_readaddr,
        doutb     => AS_D5PHIBn1_V_dout,
        sync_nent => AS_D5PHIBn1_start,
        nent_o    => AS_D5PHIBn1_AV_dout_nent
      );

    AS_D5PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIBn1_wea,
        addra     => AS_D5PHIBn1_writeaddr,
        dina      => AS_D5PHIBn1_din,
        wea_out       => AS_D5PHIBn1_wea_delay,
        addra_out     => AS_D5PHIBn1_writeaddr_delay,
        dina_out      => AS_D5PHIBn1_din_delay,
        done       => VMR_done,
        start      => AS_D5PHIBn1_start
      );

    AS_D5PHICn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D5PHICn1_bx,
        bx_vld => AS_D5PHICn1_bx_vld
      );

--    STREAM_AS_D5PHICn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D5PHICn1_bx,
--        bx_in_vld => AS_D5PHICn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D5PHICn1_stream_V_dout,
--        din0=>AS_D5PHICn1_V_dout,
--        din1=>AS_D5PHICn1_V_dout,
--        din2=>AS_D5PHICn1_V_dout,
--        din3=>AS_D5PHICn1_V_dout,
--        nent0=>AS_D5PHICn1_AV_dout_nent,
--        nent1=>AS_D5PHICn1_AV_dout_nent,
--        nent2=>AS_D5PHICn1_AV_dout_nent,
--        nent3=>AS_D5PHICn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D5PHICn1_V_readaddr
--      );

    AS_D5PHICn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHICn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHICn1_wea_delay,
        addra     => AS_D5PHICn1_writeaddr_delay,
        dina      => AS_D5PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHICn1_V_readaddr,
        doutb     => AS_D5PHICn1_V_dout,
        sync_nent => AS_D5PHICn1_start,
        nent_o    => AS_D5PHICn1_AV_dout_nent
      );

    AS_D5PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHICn1_wea,
        addra     => AS_D5PHICn1_writeaddr,
        dina      => AS_D5PHICn1_din,
        wea_out       => AS_D5PHICn1_wea_delay,
        addra_out     => AS_D5PHICn1_writeaddr_delay,
        dina_out      => AS_D5PHICn1_din_delay,
        done       => VMR_done,
        start      => AS_D5PHICn1_start
      );

    AS_D5PHIDn1_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => AS_D5PHIDn1_bx,
        bx_vld => AS_D5PHIDn1_bx_vld
      );

--    STREAM_AS_D5PHIDn1 : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 36,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 0
--      )
--      port map (
--        bx_in => AS_D5PHIDn1_bx,
--        bx_in_vld => AS_D5PHIDn1_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => AS_D5PHIDn1_stream_V_dout,
--        din0=>AS_D5PHIDn1_V_dout,
--        din1=>AS_D5PHIDn1_V_dout,
--        din2=>AS_D5PHIDn1_V_dout,
--        din3=>AS_D5PHIDn1_V_dout,
--        nent0=>AS_D5PHIDn1_AV_dout_nent,
--        nent1=>AS_D5PHIDn1_AV_dout_nent,
--        nent2=>AS_D5PHIDn1_AV_dout_nent,
--        nent3=>AS_D5PHIDn1_AV_dout_nent,
--        addr_arr(9 downto 0)=>AS_D5PHIDn1_V_readaddr
--      );

    AS_D5PHIDn1 : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D5PHIDn1"
      )
      port map (
        clka      => clk,
        wea       => AS_D5PHIDn1_wea_delay,
        addra     => AS_D5PHIDn1_writeaddr_delay,
        dina      => AS_D5PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D5PHIDn1_V_readaddr,
        doutb     => AS_D5PHIDn1_V_dout,
        sync_nent => AS_D5PHIDn1_start,
        nent_o    => AS_D5PHIDn1_AV_dout_nent
      );

    AS_D5PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D5PHIDn1_wea,
        addra     => AS_D5PHIDn1_writeaddr,
        dina      => AS_D5PHIDn1_din,
        wea_out       => AS_D5PHIDn1_wea_delay,
        addra_out     => AS_D5PHIDn1_writeaddr_delay,
        dina_out      => AS_D5PHIDn1_din_delay,
        done       => VMR_done,
        start      => AS_D5PHIDn1_start
      );

    AS_L2PHIA_B_L1A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIA_B_L1A"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIA_B_L1A_wea_delay,
        addra     => AS_L2PHIA_B_L1A_writeaddr_delay,
        dina      => AS_L2PHIA_B_L1A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIA_B_L1A_V_readaddr,
        doutb     => AS_L2PHIA_B_L1A_V_dout,
        sync_nent => AS_L2PHIA_B_L1A_start,
        nent_o    => open
      );

    AS_L2PHIA_B_L1A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIA_B_L1A_wea,
        addra     => AS_L2PHIA_B_L1A_writeaddr,
        dina      => AS_L2PHIA_B_L1A_din,
        wea_out       => AS_L2PHIA_B_L1A_wea_delay,
        addra_out     => AS_L2PHIA_B_L1A_writeaddr_delay,
        dina_out      => AS_L2PHIA_B_L1A_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIA_B_L1A_start
      );

    AS_L2PHIA_B_L1B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIA_B_L1B"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIA_B_L1B_wea_delay,
        addra     => AS_L2PHIA_B_L1B_writeaddr_delay,
        dina      => AS_L2PHIA_B_L1B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIA_B_L1B_V_readaddr,
        doutb     => AS_L2PHIA_B_L1B_V_dout,
        sync_nent => AS_L2PHIA_B_L1B_start,
        nent_o    => open
      );

    AS_L2PHIA_B_L1B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIA_B_L1B_wea,
        addra     => AS_L2PHIA_B_L1B_writeaddr,
        dina      => AS_L2PHIA_B_L1B_din,
        wea_out       => AS_L2PHIA_B_L1B_wea_delay,
        addra_out     => AS_L2PHIA_B_L1B_writeaddr_delay,
        dina_out      => AS_L2PHIA_B_L1B_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIA_B_L1B_start
      );

    AS_L2PHIA_B_L1C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIA_B_L1C"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIA_B_L1C_wea_delay,
        addra     => AS_L2PHIA_B_L1C_writeaddr_delay,
        dina      => AS_L2PHIA_B_L1C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIA_B_L1C_V_readaddr,
        doutb     => AS_L2PHIA_B_L1C_V_dout,
        sync_nent => AS_L2PHIA_B_L1C_start,
        nent_o    => open
      );

    AS_L2PHIA_B_L1C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIA_B_L1C_wea,
        addra     => AS_L2PHIA_B_L1C_writeaddr,
        dina      => AS_L2PHIA_B_L1C_din,
        wea_out       => AS_L2PHIA_B_L1C_wea_delay,
        addra_out     => AS_L2PHIA_B_L1C_writeaddr_delay,
        dina_out      => AS_L2PHIA_B_L1C_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIA_B_L1C_start
      );

    AS_L2PHIB_B_L1D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIB_B_L1D"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIB_B_L1D_wea_delay,
        addra     => AS_L2PHIB_B_L1D_writeaddr_delay,
        dina      => AS_L2PHIB_B_L1D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIB_B_L1D_V_readaddr,
        doutb     => AS_L2PHIB_B_L1D_V_dout,
        sync_nent => AS_L2PHIB_B_L1D_start,
        nent_o    => open
      );

    AS_L2PHIB_B_L1D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIB_B_L1D_wea,
        addra     => AS_L2PHIB_B_L1D_writeaddr,
        dina      => AS_L2PHIB_B_L1D_din,
        wea_out       => AS_L2PHIB_B_L1D_wea_delay,
        addra_out     => AS_L2PHIB_B_L1D_writeaddr_delay,
        dina_out      => AS_L2PHIB_B_L1D_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIB_B_L1D_start
      );

    AS_L2PHIB_B_L1E : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIB_B_L1E"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIB_B_L1E_wea_delay,
        addra     => AS_L2PHIB_B_L1E_writeaddr_delay,
        dina      => AS_L2PHIB_B_L1E_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIB_B_L1E_V_readaddr,
        doutb     => AS_L2PHIB_B_L1E_V_dout,
        sync_nent => AS_L2PHIB_B_L1E_start,
        nent_o    => open
      );

    AS_L2PHIB_B_L1E_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIB_B_L1E_wea,
        addra     => AS_L2PHIB_B_L1E_writeaddr,
        dina      => AS_L2PHIB_B_L1E_din,
        wea_out       => AS_L2PHIB_B_L1E_wea_delay,
        addra_out     => AS_L2PHIB_B_L1E_writeaddr_delay,
        dina_out      => AS_L2PHIB_B_L1E_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIB_B_L1E_start
      );

    AS_L2PHIB_B_L1F : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIB_B_L1F"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIB_B_L1F_wea_delay,
        addra     => AS_L2PHIB_B_L1F_writeaddr_delay,
        dina      => AS_L2PHIB_B_L1F_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIB_B_L1F_V_readaddr,
        doutb     => AS_L2PHIB_B_L1F_V_dout,
        sync_nent => AS_L2PHIB_B_L1F_start,
        nent_o    => open
      );

    AS_L2PHIB_B_L1F_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIB_B_L1F_wea,
        addra     => AS_L2PHIB_B_L1F_writeaddr,
        dina      => AS_L2PHIB_B_L1F_din,
        wea_out       => AS_L2PHIB_B_L1F_wea_delay,
        addra_out     => AS_L2PHIB_B_L1F_writeaddr_delay,
        dina_out      => AS_L2PHIB_B_L1F_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIB_B_L1F_start
      );

    AS_L2PHIC_B_L1G : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIC_B_L1G"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIC_B_L1G_wea_delay,
        addra     => AS_L2PHIC_B_L1G_writeaddr_delay,
        dina      => AS_L2PHIC_B_L1G_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIC_B_L1G_V_readaddr,
        doutb     => AS_L2PHIC_B_L1G_V_dout,
        sync_nent => AS_L2PHIC_B_L1G_start,
        nent_o    => open
      );

    AS_L2PHIC_B_L1G_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIC_B_L1G_wea,
        addra     => AS_L2PHIC_B_L1G_writeaddr,
        dina      => AS_L2PHIC_B_L1G_din,
        wea_out       => AS_L2PHIC_B_L1G_wea_delay,
        addra_out     => AS_L2PHIC_B_L1G_writeaddr_delay,
        dina_out      => AS_L2PHIC_B_L1G_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIC_B_L1G_start
      );

    AS_L2PHIC_B_L1H : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIC_B_L1H"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIC_B_L1H_wea_delay,
        addra     => AS_L2PHIC_B_L1H_writeaddr_delay,
        dina      => AS_L2PHIC_B_L1H_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIC_B_L1H_V_readaddr,
        doutb     => AS_L2PHIC_B_L1H_V_dout,
        sync_nent => AS_L2PHIC_B_L1H_start,
        nent_o    => open
      );

    AS_L2PHIC_B_L1H_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIC_B_L1H_wea,
        addra     => AS_L2PHIC_B_L1H_writeaddr,
        dina      => AS_L2PHIC_B_L1H_din,
        wea_out       => AS_L2PHIC_B_L1H_wea_delay,
        addra_out     => AS_L2PHIC_B_L1H_writeaddr_delay,
        dina_out      => AS_L2PHIC_B_L1H_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIC_B_L1H_start
      );

    AS_L2PHIC_B_L1I : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIC_B_L1I"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIC_B_L1I_wea_delay,
        addra     => AS_L2PHIC_B_L1I_writeaddr_delay,
        dina      => AS_L2PHIC_B_L1I_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIC_B_L1I_V_readaddr,
        doutb     => AS_L2PHIC_B_L1I_V_dout,
        sync_nent => AS_L2PHIC_B_L1I_start,
        nent_o    => open
      );

    AS_L2PHIC_B_L1I_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIC_B_L1I_wea,
        addra     => AS_L2PHIC_B_L1I_writeaddr,
        dina      => AS_L2PHIC_B_L1I_din,
        wea_out       => AS_L2PHIC_B_L1I_wea_delay,
        addra_out     => AS_L2PHIC_B_L1I_writeaddr_delay,
        dina_out      => AS_L2PHIC_B_L1I_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIC_B_L1I_start
      );

    AS_L2PHID_B_L1J : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHID_B_L1J"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHID_B_L1J_wea_delay,
        addra     => AS_L2PHID_B_L1J_writeaddr_delay,
        dina      => AS_L2PHID_B_L1J_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHID_B_L1J_V_readaddr,
        doutb     => AS_L2PHID_B_L1J_V_dout,
        sync_nent => AS_L2PHID_B_L1J_start,
        nent_o    => open
      );

    AS_L2PHID_B_L1J_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHID_B_L1J_wea,
        addra     => AS_L2PHID_B_L1J_writeaddr,
        dina      => AS_L2PHID_B_L1J_din,
        wea_out       => AS_L2PHID_B_L1J_wea_delay,
        addra_out     => AS_L2PHID_B_L1J_writeaddr_delay,
        dina_out      => AS_L2PHID_B_L1J_din_delay,
        done       => VMR_done,
        start      => AS_L2PHID_B_L1J_start
      );

    AS_L2PHID_B_L1K : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHID_B_L1K"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHID_B_L1K_wea_delay,
        addra     => AS_L2PHID_B_L1K_writeaddr_delay,
        dina      => AS_L2PHID_B_L1K_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHID_B_L1K_V_readaddr,
        doutb     => AS_L2PHID_B_L1K_V_dout,
        sync_nent => AS_L2PHID_B_L1K_start,
        nent_o    => open
      );

    AS_L2PHID_B_L1K_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHID_B_L1K_wea,
        addra     => AS_L2PHID_B_L1K_writeaddr,
        dina      => AS_L2PHID_B_L1K_din,
        wea_out       => AS_L2PHID_B_L1K_wea_delay,
        addra_out     => AS_L2PHID_B_L1K_writeaddr_delay,
        dina_out      => AS_L2PHID_B_L1K_din_delay,
        done       => VMR_done,
        start      => AS_L2PHID_B_L1K_start
      );

    AS_L2PHID_B_L1L : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHID_B_L1L"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHID_B_L1L_wea_delay,
        addra     => AS_L2PHID_B_L1L_writeaddr_delay,
        dina      => AS_L2PHID_B_L1L_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHID_B_L1L_V_readaddr,
        doutb     => AS_L2PHID_B_L1L_V_dout,
        sync_nent => AS_L2PHID_B_L1L_start,
        nent_o    => open
      );

    AS_L2PHID_B_L1L_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHID_B_L1L_wea,
        addra     => AS_L2PHID_B_L1L_writeaddr,
        dina      => AS_L2PHID_B_L1L_din,
        wea_out       => AS_L2PHID_B_L1L_wea_delay,
        addra_out     => AS_L2PHID_B_L1L_writeaddr_delay,
        dina_out      => AS_L2PHID_B_L1L_din_delay,
        done       => VMR_done,
        start      => AS_L2PHID_B_L1L_start
      );

    AS_L3PHIA_B_L2A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIA_B_L2A"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIA_B_L2A_wea_delay,
        addra     => AS_L3PHIA_B_L2A_writeaddr_delay,
        dina      => AS_L3PHIA_B_L2A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIA_B_L2A_V_readaddr,
        doutb     => AS_L3PHIA_B_L2A_V_dout,
        sync_nent => AS_L3PHIA_B_L2A_start,
        nent_o    => open
      );

    AS_L3PHIA_B_L2A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIA_B_L2A_wea,
        addra     => AS_L3PHIA_B_L2A_writeaddr,
        dina      => AS_L3PHIA_B_L2A_din,
        wea_out       => AS_L3PHIA_B_L2A_wea_delay,
        addra_out     => AS_L3PHIA_B_L2A_writeaddr_delay,
        dina_out      => AS_L3PHIA_B_L2A_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIA_B_L2A_start
      );

    AS_L3PHIB_B_L2B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIB_B_L2B"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIB_B_L2B_wea_delay,
        addra     => AS_L3PHIB_B_L2B_writeaddr_delay,
        dina      => AS_L3PHIB_B_L2B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIB_B_L2B_V_readaddr,
        doutb     => AS_L3PHIB_B_L2B_V_dout,
        sync_nent => AS_L3PHIB_B_L2B_start,
        nent_o    => open
      );

    AS_L3PHIB_B_L2B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIB_B_L2B_wea,
        addra     => AS_L3PHIB_B_L2B_writeaddr,
        dina      => AS_L3PHIB_B_L2B_din,
        wea_out       => AS_L3PHIB_B_L2B_wea_delay,
        addra_out     => AS_L3PHIB_B_L2B_writeaddr_delay,
        dina_out      => AS_L3PHIB_B_L2B_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIB_B_L2B_start
      );

    AS_L3PHIC_B_L2C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIC_B_L2C"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIC_B_L2C_wea_delay,
        addra     => AS_L3PHIC_B_L2C_writeaddr_delay,
        dina      => AS_L3PHIC_B_L2C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIC_B_L2C_V_readaddr,
        doutb     => AS_L3PHIC_B_L2C_V_dout,
        sync_nent => AS_L3PHIC_B_L2C_start,
        nent_o    => open
      );

    AS_L3PHIC_B_L2C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIC_B_L2C_wea,
        addra     => AS_L3PHIC_B_L2C_writeaddr,
        dina      => AS_L3PHIC_B_L2C_din,
        wea_out       => AS_L3PHIC_B_L2C_wea_delay,
        addra_out     => AS_L3PHIC_B_L2C_writeaddr_delay,
        dina_out      => AS_L3PHIC_B_L2C_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIC_B_L2C_start
      );

    AS_L3PHID_B_L2D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHID_B_L2D"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHID_B_L2D_wea_delay,
        addra     => AS_L3PHID_B_L2D_writeaddr_delay,
        dina      => AS_L3PHID_B_L2D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHID_B_L2D_V_readaddr,
        doutb     => AS_L3PHID_B_L2D_V_dout,
        sync_nent => AS_L3PHID_B_L2D_start,
        nent_o    => open
      );

    AS_L3PHID_B_L2D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHID_B_L2D_wea,
        addra     => AS_L3PHID_B_L2D_writeaddr,
        dina      => AS_L3PHID_B_L2D_din,
        wea_out       => AS_L3PHID_B_L2D_wea_delay,
        addra_out     => AS_L3PHID_B_L2D_writeaddr_delay,
        dina_out      => AS_L3PHID_B_L2D_din_delay,
        done       => VMR_done,
        start      => AS_L3PHID_B_L2D_start
      );

    AS_L4PHIA_B_L3A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIA_B_L3A"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIA_B_L3A_wea_delay,
        addra     => AS_L4PHIA_B_L3A_writeaddr_delay,
        dina      => AS_L4PHIA_B_L3A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIA_B_L3A_V_readaddr,
        doutb     => AS_L4PHIA_B_L3A_V_dout,
        sync_nent => AS_L4PHIA_B_L3A_start,
        nent_o    => open
      );

    AS_L4PHIA_B_L3A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIA_B_L3A_wea,
        addra     => AS_L4PHIA_B_L3A_writeaddr,
        dina      => AS_L4PHIA_B_L3A_din,
        wea_out       => AS_L4PHIA_B_L3A_wea_delay,
        addra_out     => AS_L4PHIA_B_L3A_writeaddr_delay,
        dina_out      => AS_L4PHIA_B_L3A_din_delay,
        done       => VMR_done,
        start      => AS_L4PHIA_B_L3A_start
      );

    AS_L4PHIB_B_L3B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIB_B_L3B"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIB_B_L3B_wea_delay,
        addra     => AS_L4PHIB_B_L3B_writeaddr_delay,
        dina      => AS_L4PHIB_B_L3B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIB_B_L3B_V_readaddr,
        doutb     => AS_L4PHIB_B_L3B_V_dout,
        sync_nent => AS_L4PHIB_B_L3B_start,
        nent_o    => open
      );

    AS_L4PHIB_B_L3B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIB_B_L3B_wea,
        addra     => AS_L4PHIB_B_L3B_writeaddr,
        dina      => AS_L4PHIB_B_L3B_din,
        wea_out       => AS_L4PHIB_B_L3B_wea_delay,
        addra_out     => AS_L4PHIB_B_L3B_writeaddr_delay,
        dina_out      => AS_L4PHIB_B_L3B_din_delay,
        done       => VMR_done,
        start      => AS_L4PHIB_B_L3B_start
      );

    AS_L4PHIC_B_L3C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHIC_B_L3C"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHIC_B_L3C_wea_delay,
        addra     => AS_L4PHIC_B_L3C_writeaddr_delay,
        dina      => AS_L4PHIC_B_L3C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHIC_B_L3C_V_readaddr,
        doutb     => AS_L4PHIC_B_L3C_V_dout,
        sync_nent => AS_L4PHIC_B_L3C_start,
        nent_o    => open
      );

    AS_L4PHIC_B_L3C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHIC_B_L3C_wea,
        addra     => AS_L4PHIC_B_L3C_writeaddr,
        dina      => AS_L4PHIC_B_L3C_din,
        wea_out       => AS_L4PHIC_B_L3C_wea_delay,
        addra_out     => AS_L4PHIC_B_L3C_writeaddr_delay,
        dina_out      => AS_L4PHIC_B_L3C_din_delay,
        done       => VMR_done,
        start      => AS_L4PHIC_B_L3C_start
      );

    AS_L4PHID_B_L3D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L4PHID_B_L3D"
      )
      port map (
        clka      => clk,
        wea       => AS_L4PHID_B_L3D_wea_delay,
        addra     => AS_L4PHID_B_L3D_writeaddr_delay,
        dina      => AS_L4PHID_B_L3D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L4PHID_B_L3D_V_readaddr,
        doutb     => AS_L4PHID_B_L3D_V_dout,
        sync_nent => AS_L4PHID_B_L3D_start,
        nent_o    => open
      );

    AS_L4PHID_B_L3D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L4PHID_B_L3D_wea,
        addra     => AS_L4PHID_B_L3D_writeaddr,
        dina      => AS_L4PHID_B_L3D_din,
        wea_out       => AS_L4PHID_B_L3D_wea_delay,
        addra_out     => AS_L4PHID_B_L3D_writeaddr_delay,
        dina_out      => AS_L4PHID_B_L3D_din_delay,
        done       => VMR_done,
        start      => AS_L4PHID_B_L3D_start
      );

    AS_L6PHIA_B_L5A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIA_B_L5A"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIA_B_L5A_wea_delay,
        addra     => AS_L6PHIA_B_L5A_writeaddr_delay,
        dina      => AS_L6PHIA_B_L5A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIA_B_L5A_V_readaddr,
        doutb     => AS_L6PHIA_B_L5A_V_dout,
        sync_nent => AS_L6PHIA_B_L5A_start,
        nent_o    => open
      );

    AS_L6PHIA_B_L5A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIA_B_L5A_wea,
        addra     => AS_L6PHIA_B_L5A_writeaddr,
        dina      => AS_L6PHIA_B_L5A_din,
        wea_out       => AS_L6PHIA_B_L5A_wea_delay,
        addra_out     => AS_L6PHIA_B_L5A_writeaddr_delay,
        dina_out      => AS_L6PHIA_B_L5A_din_delay,
        done       => VMR_done,
        start      => AS_L6PHIA_B_L5A_start
      );

    AS_L6PHIB_B_L5B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIB_B_L5B"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIB_B_L5B_wea_delay,
        addra     => AS_L6PHIB_B_L5B_writeaddr_delay,
        dina      => AS_L6PHIB_B_L5B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIB_B_L5B_V_readaddr,
        doutb     => AS_L6PHIB_B_L5B_V_dout,
        sync_nent => AS_L6PHIB_B_L5B_start,
        nent_o    => open
      );

    AS_L6PHIB_B_L5B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIB_B_L5B_wea,
        addra     => AS_L6PHIB_B_L5B_writeaddr,
        dina      => AS_L6PHIB_B_L5B_din,
        wea_out       => AS_L6PHIB_B_L5B_wea_delay,
        addra_out     => AS_L6PHIB_B_L5B_writeaddr_delay,
        dina_out      => AS_L6PHIB_B_L5B_din_delay,
        done       => VMR_done,
        start      => AS_L6PHIB_B_L5B_start
      );

    AS_L6PHIC_B_L5C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHIC_B_L5C"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHIC_B_L5C_wea_delay,
        addra     => AS_L6PHIC_B_L5C_writeaddr_delay,
        dina      => AS_L6PHIC_B_L5C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHIC_B_L5C_V_readaddr,
        doutb     => AS_L6PHIC_B_L5C_V_dout,
        sync_nent => AS_L6PHIC_B_L5C_start,
        nent_o    => open
      );

    AS_L6PHIC_B_L5C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHIC_B_L5C_wea,
        addra     => AS_L6PHIC_B_L5C_writeaddr,
        dina      => AS_L6PHIC_B_L5C_din,
        wea_out       => AS_L6PHIC_B_L5C_wea_delay,
        addra_out     => AS_L6PHIC_B_L5C_writeaddr_delay,
        dina_out      => AS_L6PHIC_B_L5C_din_delay,
        done       => VMR_done,
        start      => AS_L6PHIC_B_L5C_start
      );

    AS_L6PHID_B_L5D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L6PHID_B_L5D"
      )
      port map (
        clka      => clk,
        wea       => AS_L6PHID_B_L5D_wea_delay,
        addra     => AS_L6PHID_B_L5D_writeaddr_delay,
        dina      => AS_L6PHID_B_L5D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L6PHID_B_L5D_V_readaddr,
        doutb     => AS_L6PHID_B_L5D_V_dout,
        sync_nent => AS_L6PHID_B_L5D_start,
        nent_o    => open
      );

    AS_L6PHID_B_L5D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_L6PHID_B_L5D_wea,
        addra     => AS_L6PHID_B_L5D_writeaddr,
        dina      => AS_L6PHID_B_L5D_din,
        wea_out       => AS_L6PHID_B_L5D_wea_delay,
        addra_out     => AS_L6PHID_B_L5D_writeaddr_delay,
        dina_out      => AS_L6PHID_B_L5D_din_delay,
        done       => VMR_done,
        start      => AS_L6PHID_B_L5D_start
      );

    AS_D1PHIA_O_L1A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIA_O_L1A"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIA_O_L1A_wea_delay,
        addra     => AS_D1PHIA_O_L1A_writeaddr_delay,
        dina      => AS_D1PHIA_O_L1A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIA_O_L1A_V_readaddr,
        doutb     => AS_D1PHIA_O_L1A_V_dout,
        sync_nent => AS_D1PHIA_O_L1A_start,
        nent_o    => open
      );

    AS_D1PHIA_O_L1A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIA_O_L1A_wea,
        addra     => AS_D1PHIA_O_L1A_writeaddr,
        dina      => AS_D1PHIA_O_L1A_din,
        wea_out       => AS_D1PHIA_O_L1A_wea_delay,
        addra_out     => AS_D1PHIA_O_L1A_writeaddr_delay,
        dina_out      => AS_D1PHIA_O_L1A_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIA_O_L1A_start
      );

    AS_D1PHIA_O_L1B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIA_O_L1B"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIA_O_L1B_wea_delay,
        addra     => AS_D1PHIA_O_L1B_writeaddr_delay,
        dina      => AS_D1PHIA_O_L1B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIA_O_L1B_V_readaddr,
        doutb     => AS_D1PHIA_O_L1B_V_dout,
        sync_nent => AS_D1PHIA_O_L1B_start,
        nent_o    => open
      );

    AS_D1PHIA_O_L1B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIA_O_L1B_wea,
        addra     => AS_D1PHIA_O_L1B_writeaddr,
        dina      => AS_D1PHIA_O_L1B_din,
        wea_out       => AS_D1PHIA_O_L1B_wea_delay,
        addra_out     => AS_D1PHIA_O_L1B_writeaddr_delay,
        dina_out      => AS_D1PHIA_O_L1B_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIA_O_L1B_start
      );

    AS_D1PHIA_O_L2A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIA_O_L2A"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIA_O_L2A_wea_delay,
        addra     => AS_D1PHIA_O_L2A_writeaddr_delay,
        dina      => AS_D1PHIA_O_L2A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIA_O_L2A_V_readaddr,
        doutb     => AS_D1PHIA_O_L2A_V_dout,
        sync_nent => AS_D1PHIA_O_L2A_start,
        nent_o    => open
      );

    AS_D1PHIA_O_L2A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIA_O_L2A_wea,
        addra     => AS_D1PHIA_O_L2A_writeaddr,
        dina      => AS_D1PHIA_O_L2A_din,
        wea_out       => AS_D1PHIA_O_L2A_wea_delay,
        addra_out     => AS_D1PHIA_O_L2A_writeaddr_delay,
        dina_out      => AS_D1PHIA_O_L2A_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIA_O_L2A_start
      );

    AS_D1PHIB_O_L1C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIB_O_L1C"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIB_O_L1C_wea_delay,
        addra     => AS_D1PHIB_O_L1C_writeaddr_delay,
        dina      => AS_D1PHIB_O_L1C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIB_O_L1C_V_readaddr,
        doutb     => AS_D1PHIB_O_L1C_V_dout,
        sync_nent => AS_D1PHIB_O_L1C_start,
        nent_o    => open
      );

    AS_D1PHIB_O_L1C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIB_O_L1C_wea,
        addra     => AS_D1PHIB_O_L1C_writeaddr,
        dina      => AS_D1PHIB_O_L1C_din,
        wea_out       => AS_D1PHIB_O_L1C_wea_delay,
        addra_out     => AS_D1PHIB_O_L1C_writeaddr_delay,
        dina_out      => AS_D1PHIB_O_L1C_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIB_O_L1C_start
      );

    AS_D1PHIB_O_L1D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIB_O_L1D"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIB_O_L1D_wea_delay,
        addra     => AS_D1PHIB_O_L1D_writeaddr_delay,
        dina      => AS_D1PHIB_O_L1D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIB_O_L1D_V_readaddr,
        doutb     => AS_D1PHIB_O_L1D_V_dout,
        sync_nent => AS_D1PHIB_O_L1D_start,
        nent_o    => open
      );

    AS_D1PHIB_O_L1D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIB_O_L1D_wea,
        addra     => AS_D1PHIB_O_L1D_writeaddr,
        dina      => AS_D1PHIB_O_L1D_din,
        wea_out       => AS_D1PHIB_O_L1D_wea_delay,
        addra_out     => AS_D1PHIB_O_L1D_writeaddr_delay,
        dina_out      => AS_D1PHIB_O_L1D_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIB_O_L1D_start
      );

    AS_D1PHIB_O_L2B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIB_O_L2B"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIB_O_L2B_wea_delay,
        addra     => AS_D1PHIB_O_L2B_writeaddr_delay,
        dina      => AS_D1PHIB_O_L2B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIB_O_L2B_V_readaddr,
        doutb     => AS_D1PHIB_O_L2B_V_dout,
        sync_nent => AS_D1PHIB_O_L2B_start,
        nent_o    => open
      );

    AS_D1PHIB_O_L2B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIB_O_L2B_wea,
        addra     => AS_D1PHIB_O_L2B_writeaddr,
        dina      => AS_D1PHIB_O_L2B_din,
        wea_out       => AS_D1PHIB_O_L2B_wea_delay,
        addra_out     => AS_D1PHIB_O_L2B_writeaddr_delay,
        dina_out      => AS_D1PHIB_O_L2B_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIB_O_L2B_start
      );

    AS_D1PHIC_O_L1E : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIC_O_L1E"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIC_O_L1E_wea_delay,
        addra     => AS_D1PHIC_O_L1E_writeaddr_delay,
        dina      => AS_D1PHIC_O_L1E_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIC_O_L1E_V_readaddr,
        doutb     => AS_D1PHIC_O_L1E_V_dout,
        sync_nent => AS_D1PHIC_O_L1E_start,
        nent_o    => open
      );

    AS_D1PHIC_O_L1E_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIC_O_L1E_wea,
        addra     => AS_D1PHIC_O_L1E_writeaddr,
        dina      => AS_D1PHIC_O_L1E_din,
        wea_out       => AS_D1PHIC_O_L1E_wea_delay,
        addra_out     => AS_D1PHIC_O_L1E_writeaddr_delay,
        dina_out      => AS_D1PHIC_O_L1E_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIC_O_L1E_start
      );

    AS_D1PHIC_O_L1F : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIC_O_L1F"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIC_O_L1F_wea_delay,
        addra     => AS_D1PHIC_O_L1F_writeaddr_delay,
        dina      => AS_D1PHIC_O_L1F_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIC_O_L1F_V_readaddr,
        doutb     => AS_D1PHIC_O_L1F_V_dout,
        sync_nent => AS_D1PHIC_O_L1F_start,
        nent_o    => open
      );

    AS_D1PHIC_O_L1F_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIC_O_L1F_wea,
        addra     => AS_D1PHIC_O_L1F_writeaddr,
        dina      => AS_D1PHIC_O_L1F_din,
        wea_out       => AS_D1PHIC_O_L1F_wea_delay,
        addra_out     => AS_D1PHIC_O_L1F_writeaddr_delay,
        dina_out      => AS_D1PHIC_O_L1F_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIC_O_L1F_start
      );

    AS_D1PHIC_O_L2C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIC_O_L2C"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIC_O_L2C_wea_delay,
        addra     => AS_D1PHIC_O_L2C_writeaddr_delay,
        dina      => AS_D1PHIC_O_L2C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIC_O_L2C_V_readaddr,
        doutb     => AS_D1PHIC_O_L2C_V_dout,
        sync_nent => AS_D1PHIC_O_L2C_start,
        nent_o    => open
      );

    AS_D1PHIC_O_L2C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIC_O_L2C_wea,
        addra     => AS_D1PHIC_O_L2C_writeaddr,
        dina      => AS_D1PHIC_O_L2C_din,
        wea_out       => AS_D1PHIC_O_L2C_wea_delay,
        addra_out     => AS_D1PHIC_O_L2C_writeaddr_delay,
        dina_out      => AS_D1PHIC_O_L2C_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIC_O_L2C_start
      );

    AS_D1PHID_O_L1G : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHID_O_L1G"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHID_O_L1G_wea_delay,
        addra     => AS_D1PHID_O_L1G_writeaddr_delay,
        dina      => AS_D1PHID_O_L1G_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHID_O_L1G_V_readaddr,
        doutb     => AS_D1PHID_O_L1G_V_dout,
        sync_nent => AS_D1PHID_O_L1G_start,
        nent_o    => open
      );

    AS_D1PHID_O_L1G_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHID_O_L1G_wea,
        addra     => AS_D1PHID_O_L1G_writeaddr,
        dina      => AS_D1PHID_O_L1G_din,
        wea_out       => AS_D1PHID_O_L1G_wea_delay,
        addra_out     => AS_D1PHID_O_L1G_writeaddr_delay,
        dina_out      => AS_D1PHID_O_L1G_din_delay,
        done       => VMR_done,
        start      => AS_D1PHID_O_L1G_start
      );

    AS_D1PHID_O_L1H : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHID_O_L1H"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHID_O_L1H_wea_delay,
        addra     => AS_D1PHID_O_L1H_writeaddr_delay,
        dina      => AS_D1PHID_O_L1H_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHID_O_L1H_V_readaddr,
        doutb     => AS_D1PHID_O_L1H_V_dout,
        sync_nent => AS_D1PHID_O_L1H_start,
        nent_o    => open
      );

    AS_D1PHID_O_L1H_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHID_O_L1H_wea,
        addra     => AS_D1PHID_O_L1H_writeaddr,
        dina      => AS_D1PHID_O_L1H_din,
        wea_out       => AS_D1PHID_O_L1H_wea_delay,
        addra_out     => AS_D1PHID_O_L1H_writeaddr_delay,
        dina_out      => AS_D1PHID_O_L1H_din_delay,
        done       => VMR_done,
        start      => AS_D1PHID_O_L1H_start
      );

    AS_D1PHID_O_L2D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHID_O_L2D"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHID_O_L2D_wea_delay,
        addra     => AS_D1PHID_O_L2D_writeaddr_delay,
        dina      => AS_D1PHID_O_L2D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHID_O_L2D_V_readaddr,
        doutb     => AS_D1PHID_O_L2D_V_dout,
        sync_nent => AS_D1PHID_O_L2D_start,
        nent_o    => open
      );

    AS_D1PHID_O_L2D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHID_O_L2D_wea,
        addra     => AS_D1PHID_O_L2D_writeaddr,
        dina      => AS_D1PHID_O_L2D_din,
        wea_out       => AS_D1PHID_O_L2D_wea_delay,
        addra_out     => AS_D1PHID_O_L2D_writeaddr_delay,
        dina_out      => AS_D1PHID_O_L2D_din_delay,
        done       => VMR_done,
        start      => AS_D1PHID_O_L2D_start
      );

    AS_D2PHIA_D_D1A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIA_D_D1A"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIA_D_D1A_wea_delay,
        addra     => AS_D2PHIA_D_D1A_writeaddr_delay,
        dina      => AS_D2PHIA_D_D1A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIA_D_D1A_V_readaddr,
        doutb     => AS_D2PHIA_D_D1A_V_dout,
        sync_nent => AS_D2PHIA_D_D1A_start,
        nent_o    => open
      );

    AS_D2PHIA_D_D1A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIA_D_D1A_wea,
        addra     => AS_D2PHIA_D_D1A_writeaddr,
        dina      => AS_D2PHIA_D_D1A_din,
        wea_out       => AS_D2PHIA_D_D1A_wea_delay,
        addra_out     => AS_D2PHIA_D_D1A_writeaddr_delay,
        dina_out      => AS_D2PHIA_D_D1A_din_delay,
        done       => VMR_done,
        start      => AS_D2PHIA_D_D1A_start
      );

    AS_D2PHIB_D_D1B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIB_D_D1B"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIB_D_D1B_wea_delay,
        addra     => AS_D2PHIB_D_D1B_writeaddr_delay,
        dina      => AS_D2PHIB_D_D1B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIB_D_D1B_V_readaddr,
        doutb     => AS_D2PHIB_D_D1B_V_dout,
        sync_nent => AS_D2PHIB_D_D1B_start,
        nent_o    => open
      );

    AS_D2PHIB_D_D1B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIB_D_D1B_wea,
        addra     => AS_D2PHIB_D_D1B_writeaddr,
        dina      => AS_D2PHIB_D_D1B_din,
        wea_out       => AS_D2PHIB_D_D1B_wea_delay,
        addra_out     => AS_D2PHIB_D_D1B_writeaddr_delay,
        dina_out      => AS_D2PHIB_D_D1B_din_delay,
        done       => VMR_done,
        start      => AS_D2PHIB_D_D1B_start
      );

    AS_D2PHIC_D_D1C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHIC_D_D1C"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHIC_D_D1C_wea_delay,
        addra     => AS_D2PHIC_D_D1C_writeaddr_delay,
        dina      => AS_D2PHIC_D_D1C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHIC_D_D1C_V_readaddr,
        doutb     => AS_D2PHIC_D_D1C_V_dout,
        sync_nent => AS_D2PHIC_D_D1C_start,
        nent_o    => open
      );

    AS_D2PHIC_D_D1C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHIC_D_D1C_wea,
        addra     => AS_D2PHIC_D_D1C_writeaddr,
        dina      => AS_D2PHIC_D_D1C_din,
        wea_out       => AS_D2PHIC_D_D1C_wea_delay,
        addra_out     => AS_D2PHIC_D_D1C_writeaddr_delay,
        dina_out      => AS_D2PHIC_D_D1C_din_delay,
        done       => VMR_done,
        start      => AS_D2PHIC_D_D1C_start
      );

    AS_D2PHID_D_D1D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D2PHID_D_D1D"
      )
      port map (
        clka      => clk,
        wea       => AS_D2PHID_D_D1D_wea_delay,
        addra     => AS_D2PHID_D_D1D_writeaddr_delay,
        dina      => AS_D2PHID_D_D1D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D2PHID_D_D1D_V_readaddr,
        doutb     => AS_D2PHID_D_D1D_V_dout,
        sync_nent => AS_D2PHID_D_D1D_start,
        nent_o    => open
      );

    AS_D2PHID_D_D1D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D2PHID_D_D1D_wea,
        addra     => AS_D2PHID_D_D1D_writeaddr,
        dina      => AS_D2PHID_D_D1D_din,
        wea_out       => AS_D2PHID_D_D1D_wea_delay,
        addra_out     => AS_D2PHID_D_D1D_writeaddr_delay,
        dina_out      => AS_D2PHID_D_D1D_din_delay,
        done       => VMR_done,
        start      => AS_D2PHID_D_D1D_start
      );

    AS_D4PHIA_D_D3A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIA_D_D3A"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIA_D_D3A_wea_delay,
        addra     => AS_D4PHIA_D_D3A_writeaddr_delay,
        dina      => AS_D4PHIA_D_D3A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIA_D_D3A_V_readaddr,
        doutb     => AS_D4PHIA_D_D3A_V_dout,
        sync_nent => AS_D4PHIA_D_D3A_start,
        nent_o    => open
      );

    AS_D4PHIA_D_D3A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIA_D_D3A_wea,
        addra     => AS_D4PHIA_D_D3A_writeaddr,
        dina      => AS_D4PHIA_D_D3A_din,
        wea_out       => AS_D4PHIA_D_D3A_wea_delay,
        addra_out     => AS_D4PHIA_D_D3A_writeaddr_delay,
        dina_out      => AS_D4PHIA_D_D3A_din_delay,
        done       => VMR_done,
        start      => AS_D4PHIA_D_D3A_start
      );

    AS_D4PHIB_D_D3B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIB_D_D3B"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIB_D_D3B_wea_delay,
        addra     => AS_D4PHIB_D_D3B_writeaddr_delay,
        dina      => AS_D4PHIB_D_D3B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIB_D_D3B_V_readaddr,
        doutb     => AS_D4PHIB_D_D3B_V_dout,
        sync_nent => AS_D4PHIB_D_D3B_start,
        nent_o    => open
      );

    AS_D4PHIB_D_D3B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIB_D_D3B_wea,
        addra     => AS_D4PHIB_D_D3B_writeaddr,
        dina      => AS_D4PHIB_D_D3B_din,
        wea_out       => AS_D4PHIB_D_D3B_wea_delay,
        addra_out     => AS_D4PHIB_D_D3B_writeaddr_delay,
        dina_out      => AS_D4PHIB_D_D3B_din_delay,
        done       => VMR_done,
        start      => AS_D4PHIB_D_D3B_start
      );

    AS_D4PHIC_D_D3C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHIC_D_D3C"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHIC_D_D3C_wea_delay,
        addra     => AS_D4PHIC_D_D3C_writeaddr_delay,
        dina      => AS_D4PHIC_D_D3C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHIC_D_D3C_V_readaddr,
        doutb     => AS_D4PHIC_D_D3C_V_dout,
        sync_nent => AS_D4PHIC_D_D3C_start,
        nent_o    => open
      );

    AS_D4PHIC_D_D3C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHIC_D_D3C_wea,
        addra     => AS_D4PHIC_D_D3C_writeaddr,
        dina      => AS_D4PHIC_D_D3C_din,
        wea_out       => AS_D4PHIC_D_D3C_wea_delay,
        addra_out     => AS_D4PHIC_D_D3C_writeaddr_delay,
        dina_out      => AS_D4PHIC_D_D3C_din_delay,
        done       => VMR_done,
        start      => AS_D4PHIC_D_D3C_start
      );

    AS_D4PHID_D_D3D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 36,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D4PHID_D_D3D"
      )
      port map (
        clka      => clk,
        wea       => AS_D4PHID_D_D3D_wea_delay,
        addra     => AS_D4PHID_D_D3D_writeaddr_delay,
        dina      => AS_D4PHID_D_D3D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D4PHID_D_D3D_V_readaddr,
        doutb     => AS_D4PHID_D_D3D_V_dout,
        sync_nent => AS_D4PHID_D_D3D_start,
        nent_o    => open
      );

    AS_D4PHID_D_D3D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 36
      )
      port map (
        clk      => clk,
        wea       => AS_D4PHID_D_D3D_wea,
        addra     => AS_D4PHID_D_D3D_writeaddr,
        dina      => AS_D4PHID_D_D3D_din,
        wea_out       => AS_D4PHID_D_D3D_wea_delay,
        addra_out     => AS_D4PHID_D_D3D_writeaddr_delay,
        dina_out      => AS_D4PHID_D_D3D_din_delay,
        done       => VMR_done,
        start      => AS_D4PHID_D_D3D_start
      );

    AS_L1PHIA_BF : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIA_BF"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIA_BF_wea_delay,
        addra     => AS_L1PHIA_BF_writeaddr_delay,
        dina      => AS_L1PHIA_BF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIA_BF_V_readaddr,
        doutb     => AS_L1PHIA_BF_V_dout,
        sync_nent => AS_L1PHIA_BF_start,
        nent_o    => AS_L1PHIA_BF_AV_dout_nent
      );

    AS_L1PHIA_BF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIA_BF_wea,
        addra     => AS_L1PHIA_BF_writeaddr,
        dina      => AS_L1PHIA_BF_din,
        wea_out       => AS_L1PHIA_BF_wea_delay,
        addra_out     => AS_L1PHIA_BF_writeaddr_delay,
        dina_out      => AS_L1PHIA_BF_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIA_BF_start
      );

    AS_L1PHIA_BE : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIA_BE"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIA_BE_wea_delay,
        addra     => AS_L1PHIA_BE_writeaddr_delay,
        dina      => AS_L1PHIA_BE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIA_BE_V_readaddr,
        doutb     => AS_L1PHIA_BE_V_dout,
        sync_nent => AS_L1PHIA_BE_start,
        nent_o    => AS_L1PHIA_BE_AV_dout_nent
      );

    AS_L1PHIA_BE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIA_BE_wea,
        addra     => AS_L1PHIA_BE_writeaddr,
        dina      => AS_L1PHIA_BE_din,
        wea_out       => AS_L1PHIA_BE_wea_delay,
        addra_out     => AS_L1PHIA_BE_writeaddr_delay,
        dina_out      => AS_L1PHIA_BE_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIA_BE_start
      );

    AS_L1PHIA_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIA_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIA_OM_wea_delay,
        addra     => AS_L1PHIA_OM_writeaddr_delay,
        dina      => AS_L1PHIA_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIA_OM_V_readaddr,
        doutb     => AS_L1PHIA_OM_V_dout,
        sync_nent => AS_L1PHIA_OM_start,
        nent_o    => AS_L1PHIA_OM_AV_dout_nent
      );

    AS_L1PHIA_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIA_OM_wea,
        addra     => AS_L1PHIA_OM_writeaddr,
        dina      => AS_L1PHIA_OM_din,
        wea_out       => AS_L1PHIA_OM_wea_delay,
        addra_out     => AS_L1PHIA_OM_writeaddr_delay,
        dina_out      => AS_L1PHIA_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIA_OM_start
      );

    AS_L1PHIB_BD : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIB_BD"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIB_BD_wea_delay,
        addra     => AS_L1PHIB_BD_writeaddr_delay,
        dina      => AS_L1PHIB_BD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIB_BD_V_readaddr,
        doutb     => AS_L1PHIB_BD_V_dout,
        sync_nent => AS_L1PHIB_BD_start,
        nent_o    => AS_L1PHIB_BD_AV_dout_nent
      );

    AS_L1PHIB_BD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIB_BD_wea,
        addra     => AS_L1PHIB_BD_writeaddr,
        dina      => AS_L1PHIB_BD_din,
        wea_out       => AS_L1PHIB_BD_wea_delay,
        addra_out     => AS_L1PHIB_BD_writeaddr_delay,
        dina_out      => AS_L1PHIB_BD_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIB_BD_start
      );

    AS_L1PHIB_BC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIB_BC"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIB_BC_wea_delay,
        addra     => AS_L1PHIB_BC_writeaddr_delay,
        dina      => AS_L1PHIB_BC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIB_BC_V_readaddr,
        doutb     => AS_L1PHIB_BC_V_dout,
        sync_nent => AS_L1PHIB_BC_start,
        nent_o    => AS_L1PHIB_BC_AV_dout_nent
      );

    AS_L1PHIB_BC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIB_BC_wea,
        addra     => AS_L1PHIB_BC_writeaddr,
        dina      => AS_L1PHIB_BC_din,
        wea_out       => AS_L1PHIB_BC_wea_delay,
        addra_out     => AS_L1PHIB_BC_writeaddr_delay,
        dina_out      => AS_L1PHIB_BC_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIB_BC_start
      );

    AS_L1PHIB_BA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIB_BA"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIB_BA_wea_delay,
        addra     => AS_L1PHIB_BA_writeaddr_delay,
        dina      => AS_L1PHIB_BA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIB_BA_V_readaddr,
        doutb     => AS_L1PHIB_BA_V_dout,
        sync_nent => AS_L1PHIB_BA_start,
        nent_o    => AS_L1PHIB_BA_AV_dout_nent
      );

    AS_L1PHIB_BA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIB_BA_wea,
        addra     => AS_L1PHIB_BA_writeaddr,
        dina      => AS_L1PHIB_BA_din,
        wea_out       => AS_L1PHIB_BA_wea_delay,
        addra_out     => AS_L1PHIB_BA_writeaddr_delay,
        dina_out      => AS_L1PHIB_BA_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIB_BA_start
      );

    AS_L1PHIB_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIB_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIB_OM_wea_delay,
        addra     => AS_L1PHIB_OM_writeaddr_delay,
        dina      => AS_L1PHIB_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIB_OM_V_readaddr,
        doutb     => AS_L1PHIB_OM_V_dout,
        sync_nent => AS_L1PHIB_OM_start,
        nent_o    => AS_L1PHIB_OM_AV_dout_nent
      );

    AS_L1PHIB_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIB_OM_wea,
        addra     => AS_L1PHIB_OM_writeaddr,
        dina      => AS_L1PHIB_OM_din,
        wea_out       => AS_L1PHIB_OM_wea_delay,
        addra_out     => AS_L1PHIB_OM_writeaddr_delay,
        dina_out      => AS_L1PHIB_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIB_OM_start
      );

    AS_L1PHIB_OR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIB_OR"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIB_OR_wea_delay,
        addra     => AS_L1PHIB_OR_writeaddr_delay,
        dina      => AS_L1PHIB_OR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIB_OR_V_readaddr,
        doutb     => AS_L1PHIB_OR_V_dout,
        sync_nent => AS_L1PHIB_OR_start,
        nent_o    => AS_L1PHIB_OR_AV_dout_nent
      );

    AS_L1PHIB_OR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIB_OR_wea,
        addra     => AS_L1PHIB_OR_writeaddr,
        dina      => AS_L1PHIB_OR_din,
        wea_out       => AS_L1PHIB_OR_wea_delay,
        addra_out     => AS_L1PHIB_OR_writeaddr_delay,
        dina_out      => AS_L1PHIB_OR_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIB_OR_start
      );

    AS_L1PHIC_BB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIC_BB"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIC_BB_wea_delay,
        addra     => AS_L1PHIC_BB_writeaddr_delay,
        dina      => AS_L1PHIC_BB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIC_BB_V_readaddr,
        doutb     => AS_L1PHIC_BB_V_dout,
        sync_nent => AS_L1PHIC_BB_start,
        nent_o    => AS_L1PHIC_BB_AV_dout_nent
      );

    AS_L1PHIC_BB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIC_BB_wea,
        addra     => AS_L1PHIC_BB_writeaddr,
        dina      => AS_L1PHIC_BB_din,
        wea_out       => AS_L1PHIC_BB_wea_delay,
        addra_out     => AS_L1PHIC_BB_writeaddr_delay,
        dina_out      => AS_L1PHIC_BB_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIC_BB_start
      );

    AS_L1PHIC_BF : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIC_BF"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIC_BF_wea_delay,
        addra     => AS_L1PHIC_BF_writeaddr_delay,
        dina      => AS_L1PHIC_BF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIC_BF_V_readaddr,
        doutb     => AS_L1PHIC_BF_V_dout,
        sync_nent => AS_L1PHIC_BF_start,
        nent_o    => AS_L1PHIC_BF_AV_dout_nent
      );

    AS_L1PHIC_BF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIC_BF_wea,
        addra     => AS_L1PHIC_BF_writeaddr,
        dina      => AS_L1PHIC_BF_din,
        wea_out       => AS_L1PHIC_BF_wea_delay,
        addra_out     => AS_L1PHIC_BF_writeaddr_delay,
        dina_out      => AS_L1PHIC_BF_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIC_BF_start
      );

    AS_L1PHIC_BE : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIC_BE"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIC_BE_wea_delay,
        addra     => AS_L1PHIC_BE_writeaddr_delay,
        dina      => AS_L1PHIC_BE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIC_BE_V_readaddr,
        doutb     => AS_L1PHIC_BE_V_dout,
        sync_nent => AS_L1PHIC_BE_start,
        nent_o    => AS_L1PHIC_BE_AV_dout_nent
      );

    AS_L1PHIC_BE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIC_BE_wea,
        addra     => AS_L1PHIC_BE_writeaddr,
        dina      => AS_L1PHIC_BE_din,
        wea_out       => AS_L1PHIC_BE_wea_delay,
        addra_out     => AS_L1PHIC_BE_writeaddr_delay,
        dina_out      => AS_L1PHIC_BE_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIC_BE_start
      );

    AS_L1PHIC_OL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIC_OL"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIC_OL_wea_delay,
        addra     => AS_L1PHIC_OL_writeaddr_delay,
        dina      => AS_L1PHIC_OL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIC_OL_V_readaddr,
        doutb     => AS_L1PHIC_OL_V_dout,
        sync_nent => AS_L1PHIC_OL_start,
        nent_o    => AS_L1PHIC_OL_AV_dout_nent
      );

    AS_L1PHIC_OL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIC_OL_wea,
        addra     => AS_L1PHIC_OL_writeaddr,
        dina      => AS_L1PHIC_OL_din,
        wea_out       => AS_L1PHIC_OL_wea_delay,
        addra_out     => AS_L1PHIC_OL_writeaddr_delay,
        dina_out      => AS_L1PHIC_OL_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIC_OL_start
      );

    AS_L1PHIC_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIC_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIC_OM_wea_delay,
        addra     => AS_L1PHIC_OM_writeaddr_delay,
        dina      => AS_L1PHIC_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIC_OM_V_readaddr,
        doutb     => AS_L1PHIC_OM_V_dout,
        sync_nent => AS_L1PHIC_OM_start,
        nent_o    => AS_L1PHIC_OM_AV_dout_nent
      );

    AS_L1PHIC_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIC_OM_wea,
        addra     => AS_L1PHIC_OM_writeaddr,
        dina      => AS_L1PHIC_OM_din,
        wea_out       => AS_L1PHIC_OM_wea_delay,
        addra_out     => AS_L1PHIC_OM_writeaddr_delay,
        dina_out      => AS_L1PHIC_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIC_OM_start
      );

    AS_L1PHID_BD : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHID_BD"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHID_BD_wea_delay,
        addra     => AS_L1PHID_BD_writeaddr_delay,
        dina      => AS_L1PHID_BD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHID_BD_V_readaddr,
        doutb     => AS_L1PHID_BD_V_dout,
        sync_nent => AS_L1PHID_BD_start,
        nent_o    => AS_L1PHID_BD_AV_dout_nent
      );

    AS_L1PHID_BD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHID_BD_wea,
        addra     => AS_L1PHID_BD_writeaddr,
        dina      => AS_L1PHID_BD_din,
        wea_out       => AS_L1PHID_BD_wea_delay,
        addra_out     => AS_L1PHID_BD_writeaddr_delay,
        dina_out      => AS_L1PHID_BD_din_delay,
        done       => VMR_done,
        start      => AS_L1PHID_BD_start
      );

    AS_L1PHID_BC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHID_BC"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHID_BC_wea_delay,
        addra     => AS_L1PHID_BC_writeaddr_delay,
        dina      => AS_L1PHID_BC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHID_BC_V_readaddr,
        doutb     => AS_L1PHID_BC_V_dout,
        sync_nent => AS_L1PHID_BC_start,
        nent_o    => AS_L1PHID_BC_AV_dout_nent
      );

    AS_L1PHID_BC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHID_BC_wea,
        addra     => AS_L1PHID_BC_writeaddr,
        dina      => AS_L1PHID_BC_din,
        wea_out       => AS_L1PHID_BC_wea_delay,
        addra_out     => AS_L1PHID_BC_writeaddr_delay,
        dina_out      => AS_L1PHID_BC_din_delay,
        done       => VMR_done,
        start      => AS_L1PHID_BC_start
      );

    AS_L1PHID_BA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHID_BA"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHID_BA_wea_delay,
        addra     => AS_L1PHID_BA_writeaddr_delay,
        dina      => AS_L1PHID_BA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHID_BA_V_readaddr,
        doutb     => AS_L1PHID_BA_V_dout,
        sync_nent => AS_L1PHID_BA_start,
        nent_o    => AS_L1PHID_BA_AV_dout_nent
      );

    AS_L1PHID_BA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHID_BA_wea,
        addra     => AS_L1PHID_BA_writeaddr,
        dina      => AS_L1PHID_BA_din,
        wea_out       => AS_L1PHID_BA_wea_delay,
        addra_out     => AS_L1PHID_BA_writeaddr_delay,
        dina_out      => AS_L1PHID_BA_din_delay,
        done       => VMR_done,
        start      => AS_L1PHID_BA_start
      );

    AS_L1PHID_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHID_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHID_OM_wea_delay,
        addra     => AS_L1PHID_OM_writeaddr_delay,
        dina      => AS_L1PHID_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHID_OM_V_readaddr,
        doutb     => AS_L1PHID_OM_V_dout,
        sync_nent => AS_L1PHID_OM_start,
        nent_o    => AS_L1PHID_OM_AV_dout_nent
      );

    AS_L1PHID_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHID_OM_wea,
        addra     => AS_L1PHID_OM_writeaddr,
        dina      => AS_L1PHID_OM_din,
        wea_out       => AS_L1PHID_OM_wea_delay,
        addra_out     => AS_L1PHID_OM_writeaddr_delay,
        dina_out      => AS_L1PHID_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHID_OM_start
      );

    AS_L1PHID_OR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHID_OR"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHID_OR_wea_delay,
        addra     => AS_L1PHID_OR_writeaddr_delay,
        dina      => AS_L1PHID_OR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHID_OR_V_readaddr,
        doutb     => AS_L1PHID_OR_V_dout,
        sync_nent => AS_L1PHID_OR_start,
        nent_o    => AS_L1PHID_OR_AV_dout_nent
      );

    AS_L1PHID_OR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHID_OR_wea,
        addra     => AS_L1PHID_OR_writeaddr,
        dina      => AS_L1PHID_OR_din,
        wea_out       => AS_L1PHID_OR_wea_delay,
        addra_out     => AS_L1PHID_OR_writeaddr_delay,
        dina_out      => AS_L1PHID_OR_din_delay,
        done       => VMR_done,
        start      => AS_L1PHID_OR_start
      );

    AS_L1PHIE_BB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIE_BB"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIE_BB_wea_delay,
        addra     => AS_L1PHIE_BB_writeaddr_delay,
        dina      => AS_L1PHIE_BB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIE_BB_V_readaddr,
        doutb     => AS_L1PHIE_BB_V_dout,
        sync_nent => AS_L1PHIE_BB_start,
        nent_o    => AS_L1PHIE_BB_AV_dout_nent
      );

    AS_L1PHIE_BB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIE_BB_wea,
        addra     => AS_L1PHIE_BB_writeaddr,
        dina      => AS_L1PHIE_BB_din,
        wea_out       => AS_L1PHIE_BB_wea_delay,
        addra_out     => AS_L1PHIE_BB_writeaddr_delay,
        dina_out      => AS_L1PHIE_BB_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIE_BB_start
      );

    AS_L1PHIE_BF : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIE_BF"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIE_BF_wea_delay,
        addra     => AS_L1PHIE_BF_writeaddr_delay,
        dina      => AS_L1PHIE_BF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIE_BF_V_readaddr,
        doutb     => AS_L1PHIE_BF_V_dout,
        sync_nent => AS_L1PHIE_BF_start,
        nent_o    => AS_L1PHIE_BF_AV_dout_nent
      );

    AS_L1PHIE_BF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIE_BF_wea,
        addra     => AS_L1PHIE_BF_writeaddr,
        dina      => AS_L1PHIE_BF_din,
        wea_out       => AS_L1PHIE_BF_wea_delay,
        addra_out     => AS_L1PHIE_BF_writeaddr_delay,
        dina_out      => AS_L1PHIE_BF_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIE_BF_start
      );

    AS_L1PHIE_BE : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIE_BE"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIE_BE_wea_delay,
        addra     => AS_L1PHIE_BE_writeaddr_delay,
        dina      => AS_L1PHIE_BE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIE_BE_V_readaddr,
        doutb     => AS_L1PHIE_BE_V_dout,
        sync_nent => AS_L1PHIE_BE_start,
        nent_o    => AS_L1PHIE_BE_AV_dout_nent
      );

    AS_L1PHIE_BE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIE_BE_wea,
        addra     => AS_L1PHIE_BE_writeaddr,
        dina      => AS_L1PHIE_BE_din,
        wea_out       => AS_L1PHIE_BE_wea_delay,
        addra_out     => AS_L1PHIE_BE_writeaddr_delay,
        dina_out      => AS_L1PHIE_BE_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIE_BE_start
      );

    AS_L1PHIE_OL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIE_OL"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIE_OL_wea_delay,
        addra     => AS_L1PHIE_OL_writeaddr_delay,
        dina      => AS_L1PHIE_OL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIE_OL_V_readaddr,
        doutb     => AS_L1PHIE_OL_V_dout,
        sync_nent => AS_L1PHIE_OL_start,
        nent_o    => AS_L1PHIE_OL_AV_dout_nent
      );

    AS_L1PHIE_OL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIE_OL_wea,
        addra     => AS_L1PHIE_OL_writeaddr,
        dina      => AS_L1PHIE_OL_din,
        wea_out       => AS_L1PHIE_OL_wea_delay,
        addra_out     => AS_L1PHIE_OL_writeaddr_delay,
        dina_out      => AS_L1PHIE_OL_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIE_OL_start
      );

    AS_L1PHIE_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIE_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIE_OM_wea_delay,
        addra     => AS_L1PHIE_OM_writeaddr_delay,
        dina      => AS_L1PHIE_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIE_OM_V_readaddr,
        doutb     => AS_L1PHIE_OM_V_dout,
        sync_nent => AS_L1PHIE_OM_start,
        nent_o    => AS_L1PHIE_OM_AV_dout_nent
      );

    AS_L1PHIE_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIE_OM_wea,
        addra     => AS_L1PHIE_OM_writeaddr,
        dina      => AS_L1PHIE_OM_din,
        wea_out       => AS_L1PHIE_OM_wea_delay,
        addra_out     => AS_L1PHIE_OM_writeaddr_delay,
        dina_out      => AS_L1PHIE_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIE_OM_start
      );

    AS_L1PHIF_BD : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIF_BD"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIF_BD_wea_delay,
        addra     => AS_L1PHIF_BD_writeaddr_delay,
        dina      => AS_L1PHIF_BD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIF_BD_V_readaddr,
        doutb     => AS_L1PHIF_BD_V_dout,
        sync_nent => AS_L1PHIF_BD_start,
        nent_o    => AS_L1PHIF_BD_AV_dout_nent
      );

    AS_L1PHIF_BD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIF_BD_wea,
        addra     => AS_L1PHIF_BD_writeaddr,
        dina      => AS_L1PHIF_BD_din,
        wea_out       => AS_L1PHIF_BD_wea_delay,
        addra_out     => AS_L1PHIF_BD_writeaddr_delay,
        dina_out      => AS_L1PHIF_BD_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIF_BD_start
      );

    AS_L1PHIF_BC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIF_BC"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIF_BC_wea_delay,
        addra     => AS_L1PHIF_BC_writeaddr_delay,
        dina      => AS_L1PHIF_BC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIF_BC_V_readaddr,
        doutb     => AS_L1PHIF_BC_V_dout,
        sync_nent => AS_L1PHIF_BC_start,
        nent_o    => AS_L1PHIF_BC_AV_dout_nent
      );

    AS_L1PHIF_BC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIF_BC_wea,
        addra     => AS_L1PHIF_BC_writeaddr,
        dina      => AS_L1PHIF_BC_din,
        wea_out       => AS_L1PHIF_BC_wea_delay,
        addra_out     => AS_L1PHIF_BC_writeaddr_delay,
        dina_out      => AS_L1PHIF_BC_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIF_BC_start
      );

    AS_L1PHIF_BA : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIF_BA"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIF_BA_wea_delay,
        addra     => AS_L1PHIF_BA_writeaddr_delay,
        dina      => AS_L1PHIF_BA_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIF_BA_V_readaddr,
        doutb     => AS_L1PHIF_BA_V_dout,
        sync_nent => AS_L1PHIF_BA_start,
        nent_o    => AS_L1PHIF_BA_AV_dout_nent
      );

    AS_L1PHIF_BA_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIF_BA_wea,
        addra     => AS_L1PHIF_BA_writeaddr,
        dina      => AS_L1PHIF_BA_din,
        wea_out       => AS_L1PHIF_BA_wea_delay,
        addra_out     => AS_L1PHIF_BA_writeaddr_delay,
        dina_out      => AS_L1PHIF_BA_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIF_BA_start
      );

    AS_L1PHIF_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIF_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIF_OM_wea_delay,
        addra     => AS_L1PHIF_OM_writeaddr_delay,
        dina      => AS_L1PHIF_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIF_OM_V_readaddr,
        doutb     => AS_L1PHIF_OM_V_dout,
        sync_nent => AS_L1PHIF_OM_start,
        nent_o    => AS_L1PHIF_OM_AV_dout_nent
      );

    AS_L1PHIF_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIF_OM_wea,
        addra     => AS_L1PHIF_OM_writeaddr,
        dina      => AS_L1PHIF_OM_din,
        wea_out       => AS_L1PHIF_OM_wea_delay,
        addra_out     => AS_L1PHIF_OM_writeaddr_delay,
        dina_out      => AS_L1PHIF_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIF_OM_start
      );

    AS_L1PHIF_OR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIF_OR"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIF_OR_wea_delay,
        addra     => AS_L1PHIF_OR_writeaddr_delay,
        dina      => AS_L1PHIF_OR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIF_OR_V_readaddr,
        doutb     => AS_L1PHIF_OR_V_dout,
        sync_nent => AS_L1PHIF_OR_start,
        nent_o    => AS_L1PHIF_OR_AV_dout_nent
      );

    AS_L1PHIF_OR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIF_OR_wea,
        addra     => AS_L1PHIF_OR_writeaddr,
        dina      => AS_L1PHIF_OR_din,
        wea_out       => AS_L1PHIF_OR_wea_delay,
        addra_out     => AS_L1PHIF_OR_writeaddr_delay,
        dina_out      => AS_L1PHIF_OR_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIF_OR_start
      );

    AS_L1PHIG_BB : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIG_BB"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIG_BB_wea_delay,
        addra     => AS_L1PHIG_BB_writeaddr_delay,
        dina      => AS_L1PHIG_BB_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIG_BB_V_readaddr,
        doutb     => AS_L1PHIG_BB_V_dout,
        sync_nent => AS_L1PHIG_BB_start,
        nent_o    => AS_L1PHIG_BB_AV_dout_nent
      );

    AS_L1PHIG_BB_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIG_BB_wea,
        addra     => AS_L1PHIG_BB_writeaddr,
        dina      => AS_L1PHIG_BB_din,
        wea_out       => AS_L1PHIG_BB_wea_delay,
        addra_out     => AS_L1PHIG_BB_writeaddr_delay,
        dina_out      => AS_L1PHIG_BB_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIG_BB_start
      );

    AS_L1PHIG_BF : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIG_BF"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIG_BF_wea_delay,
        addra     => AS_L1PHIG_BF_writeaddr_delay,
        dina      => AS_L1PHIG_BF_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIG_BF_V_readaddr,
        doutb     => AS_L1PHIG_BF_V_dout,
        sync_nent => AS_L1PHIG_BF_start,
        nent_o    => AS_L1PHIG_BF_AV_dout_nent
      );

    AS_L1PHIG_BF_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIG_BF_wea,
        addra     => AS_L1PHIG_BF_writeaddr,
        dina      => AS_L1PHIG_BF_din,
        wea_out       => AS_L1PHIG_BF_wea_delay,
        addra_out     => AS_L1PHIG_BF_writeaddr_delay,
        dina_out      => AS_L1PHIG_BF_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIG_BF_start
      );

    AS_L1PHIG_BE : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIG_BE"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIG_BE_wea_delay,
        addra     => AS_L1PHIG_BE_writeaddr_delay,
        dina      => AS_L1PHIG_BE_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIG_BE_V_readaddr,
        doutb     => AS_L1PHIG_BE_V_dout,
        sync_nent => AS_L1PHIG_BE_start,
        nent_o    => AS_L1PHIG_BE_AV_dout_nent
      );

    AS_L1PHIG_BE_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIG_BE_wea,
        addra     => AS_L1PHIG_BE_writeaddr,
        dina      => AS_L1PHIG_BE_din,
        wea_out       => AS_L1PHIG_BE_wea_delay,
        addra_out     => AS_L1PHIG_BE_writeaddr_delay,
        dina_out      => AS_L1PHIG_BE_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIG_BE_start
      );

    AS_L1PHIG_OL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIG_OL"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIG_OL_wea_delay,
        addra     => AS_L1PHIG_OL_writeaddr_delay,
        dina      => AS_L1PHIG_OL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIG_OL_V_readaddr,
        doutb     => AS_L1PHIG_OL_V_dout,
        sync_nent => AS_L1PHIG_OL_start,
        nent_o    => AS_L1PHIG_OL_AV_dout_nent
      );

    AS_L1PHIG_OL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIG_OL_wea,
        addra     => AS_L1PHIG_OL_writeaddr,
        dina      => AS_L1PHIG_OL_din,
        wea_out       => AS_L1PHIG_OL_wea_delay,
        addra_out     => AS_L1PHIG_OL_writeaddr_delay,
        dina_out      => AS_L1PHIG_OL_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIG_OL_start
      );

    AS_L1PHIG_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIG_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIG_OM_wea_delay,
        addra     => AS_L1PHIG_OM_writeaddr_delay,
        dina      => AS_L1PHIG_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIG_OM_V_readaddr,
        doutb     => AS_L1PHIG_OM_V_dout,
        sync_nent => AS_L1PHIG_OM_start,
        nent_o    => AS_L1PHIG_OM_AV_dout_nent
      );

    AS_L1PHIG_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIG_OM_wea,
        addra     => AS_L1PHIG_OM_writeaddr,
        dina      => AS_L1PHIG_OM_din,
        wea_out       => AS_L1PHIG_OM_wea_delay,
        addra_out     => AS_L1PHIG_OM_writeaddr_delay,
        dina_out      => AS_L1PHIG_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIG_OM_start
      );

    AS_L1PHIH_BD : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIH_BD"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIH_BD_wea_delay,
        addra     => AS_L1PHIH_BD_writeaddr_delay,
        dina      => AS_L1PHIH_BD_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIH_BD_V_readaddr,
        doutb     => AS_L1PHIH_BD_V_dout,
        sync_nent => AS_L1PHIH_BD_start,
        nent_o    => AS_L1PHIH_BD_AV_dout_nent
      );

    AS_L1PHIH_BD_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIH_BD_wea,
        addra     => AS_L1PHIH_BD_writeaddr,
        dina      => AS_L1PHIH_BD_din,
        wea_out       => AS_L1PHIH_BD_wea_delay,
        addra_out     => AS_L1PHIH_BD_writeaddr_delay,
        dina_out      => AS_L1PHIH_BD_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIH_BD_start
      );

    AS_L1PHIH_BC : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIH_BC"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIH_BC_wea_delay,
        addra     => AS_L1PHIH_BC_writeaddr_delay,
        dina      => AS_L1PHIH_BC_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIH_BC_V_readaddr,
        doutb     => AS_L1PHIH_BC_V_dout,
        sync_nent => AS_L1PHIH_BC_start,
        nent_o    => AS_L1PHIH_BC_AV_dout_nent
      );

    AS_L1PHIH_BC_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIH_BC_wea,
        addra     => AS_L1PHIH_BC_writeaddr,
        dina      => AS_L1PHIH_BC_din,
        wea_out       => AS_L1PHIH_BC_wea_delay,
        addra_out     => AS_L1PHIH_BC_writeaddr_delay,
        dina_out      => AS_L1PHIH_BC_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIH_BC_start
      );

    AS_L1PHIH_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L1PHIH_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L1PHIH_OM_wea_delay,
        addra     => AS_L1PHIH_OM_writeaddr_delay,
        dina      => AS_L1PHIH_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L1PHIH_OM_V_readaddr,
        doutb     => AS_L1PHIH_OM_V_dout,
        sync_nent => AS_L1PHIH_OM_start,
        nent_o    => AS_L1PHIH_OM_AV_dout_nent
      );

    AS_L1PHIH_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L1PHIH_OM_wea,
        addra     => AS_L1PHIH_OM_writeaddr,
        dina      => AS_L1PHIH_OM_din,
        wea_out       => AS_L1PHIH_OM_wea_delay,
        addra_out     => AS_L1PHIH_OM_writeaddr_delay,
        dina_out      => AS_L1PHIH_OM_din_delay,
        done       => VMR_done,
        start      => AS_L1PHIH_OM_start
      );

    AS_L2PHIA_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIA_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIA_BM_wea_delay,
        addra     => AS_L2PHIA_BM_writeaddr_delay,
        dina      => AS_L2PHIA_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIA_BM_V_readaddr,
        doutb     => AS_L2PHIA_BM_V_dout,
        sync_nent => AS_L2PHIA_BM_start,
        nent_o    => AS_L2PHIA_BM_AV_dout_nent
      );

    AS_L2PHIA_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIA_BM_wea,
        addra     => AS_L2PHIA_BM_writeaddr,
        dina      => AS_L2PHIA_BM_din,
        wea_out       => AS_L2PHIA_BM_wea_delay,
        addra_out     => AS_L2PHIA_BM_writeaddr_delay,
        dina_out      => AS_L2PHIA_BM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIA_BM_start
      );

    AS_L2PHIA_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIA_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIA_OM_wea_delay,
        addra     => AS_L2PHIA_OM_writeaddr_delay,
        dina      => AS_L2PHIA_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIA_OM_V_readaddr,
        doutb     => AS_L2PHIA_OM_V_dout,
        sync_nent => AS_L2PHIA_OM_start,
        nent_o    => AS_L2PHIA_OM_AV_dout_nent
      );

    AS_L2PHIA_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIA_OM_wea,
        addra     => AS_L2PHIA_OM_writeaddr,
        dina      => AS_L2PHIA_OM_din,
        wea_out       => AS_L2PHIA_OM_wea_delay,
        addra_out     => AS_L2PHIA_OM_writeaddr_delay,
        dina_out      => AS_L2PHIA_OM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIA_OM_start
      );

    AS_L2PHIB_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIB_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIB_BM_wea_delay,
        addra     => AS_L2PHIB_BM_writeaddr_delay,
        dina      => AS_L2PHIB_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIB_BM_V_readaddr,
        doutb     => AS_L2PHIB_BM_V_dout,
        sync_nent => AS_L2PHIB_BM_start,
        nent_o    => AS_L2PHIB_BM_AV_dout_nent
      );

    AS_L2PHIB_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIB_BM_wea,
        addra     => AS_L2PHIB_BM_writeaddr,
        dina      => AS_L2PHIB_BM_din,
        wea_out       => AS_L2PHIB_BM_wea_delay,
        addra_out     => AS_L2PHIB_BM_writeaddr_delay,
        dina_out      => AS_L2PHIB_BM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIB_BM_start
      );

    AS_L2PHIB_BR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIB_BR"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIB_BR_wea_delay,
        addra     => AS_L2PHIB_BR_writeaddr_delay,
        dina      => AS_L2PHIB_BR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIB_BR_V_readaddr,
        doutb     => AS_L2PHIB_BR_V_dout,
        sync_nent => AS_L2PHIB_BR_start,
        nent_o    => AS_L2PHIB_BR_AV_dout_nent
      );

    AS_L2PHIB_BR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIB_BR_wea,
        addra     => AS_L2PHIB_BR_writeaddr,
        dina      => AS_L2PHIB_BR_din,
        wea_out       => AS_L2PHIB_BR_wea_delay,
        addra_out     => AS_L2PHIB_BR_writeaddr_delay,
        dina_out      => AS_L2PHIB_BR_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIB_BR_start
      );

    AS_L2PHIB_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIB_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIB_OM_wea_delay,
        addra     => AS_L2PHIB_OM_writeaddr_delay,
        dina      => AS_L2PHIB_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIB_OM_V_readaddr,
        doutb     => AS_L2PHIB_OM_V_dout,
        sync_nent => AS_L2PHIB_OM_start,
        nent_o    => AS_L2PHIB_OM_AV_dout_nent
      );

    AS_L2PHIB_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIB_OM_wea,
        addra     => AS_L2PHIB_OM_writeaddr,
        dina      => AS_L2PHIB_OM_din,
        wea_out       => AS_L2PHIB_OM_wea_delay,
        addra_out     => AS_L2PHIB_OM_writeaddr_delay,
        dina_out      => AS_L2PHIB_OM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIB_OM_start
      );

    AS_L2PHIB_OR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIB_OR"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIB_OR_wea_delay,
        addra     => AS_L2PHIB_OR_writeaddr_delay,
        dina      => AS_L2PHIB_OR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIB_OR_V_readaddr,
        doutb     => AS_L2PHIB_OR_V_dout,
        sync_nent => AS_L2PHIB_OR_start,
        nent_o    => AS_L2PHIB_OR_AV_dout_nent
      );

    AS_L2PHIB_OR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIB_OR_wea,
        addra     => AS_L2PHIB_OR_writeaddr,
        dina      => AS_L2PHIB_OR_din,
        wea_out       => AS_L2PHIB_OR_wea_delay,
        addra_out     => AS_L2PHIB_OR_writeaddr_delay,
        dina_out      => AS_L2PHIB_OR_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIB_OR_start
      );

    AS_L2PHIC_BL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIC_BL"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIC_BL_wea_delay,
        addra     => AS_L2PHIC_BL_writeaddr_delay,
        dina      => AS_L2PHIC_BL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIC_BL_V_readaddr,
        doutb     => AS_L2PHIC_BL_V_dout,
        sync_nent => AS_L2PHIC_BL_start,
        nent_o    => AS_L2PHIC_BL_AV_dout_nent
      );

    AS_L2PHIC_BL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIC_BL_wea,
        addra     => AS_L2PHIC_BL_writeaddr,
        dina      => AS_L2PHIC_BL_din,
        wea_out       => AS_L2PHIC_BL_wea_delay,
        addra_out     => AS_L2PHIC_BL_writeaddr_delay,
        dina_out      => AS_L2PHIC_BL_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIC_BL_start
      );

    AS_L2PHIC_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIC_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIC_BM_wea_delay,
        addra     => AS_L2PHIC_BM_writeaddr_delay,
        dina      => AS_L2PHIC_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIC_BM_V_readaddr,
        doutb     => AS_L2PHIC_BM_V_dout,
        sync_nent => AS_L2PHIC_BM_start,
        nent_o    => AS_L2PHIC_BM_AV_dout_nent
      );

    AS_L2PHIC_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIC_BM_wea,
        addra     => AS_L2PHIC_BM_writeaddr,
        dina      => AS_L2PHIC_BM_din,
        wea_out       => AS_L2PHIC_BM_wea_delay,
        addra_out     => AS_L2PHIC_BM_writeaddr_delay,
        dina_out      => AS_L2PHIC_BM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIC_BM_start
      );

    AS_L2PHIC_OL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIC_OL"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIC_OL_wea_delay,
        addra     => AS_L2PHIC_OL_writeaddr_delay,
        dina      => AS_L2PHIC_OL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIC_OL_V_readaddr,
        doutb     => AS_L2PHIC_OL_V_dout,
        sync_nent => AS_L2PHIC_OL_start,
        nent_o    => AS_L2PHIC_OL_AV_dout_nent
      );

    AS_L2PHIC_OL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIC_OL_wea,
        addra     => AS_L2PHIC_OL_writeaddr,
        dina      => AS_L2PHIC_OL_din,
        wea_out       => AS_L2PHIC_OL_wea_delay,
        addra_out     => AS_L2PHIC_OL_writeaddr_delay,
        dina_out      => AS_L2PHIC_OL_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIC_OL_start
      );

    AS_L2PHIC_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHIC_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHIC_OM_wea_delay,
        addra     => AS_L2PHIC_OM_writeaddr_delay,
        dina      => AS_L2PHIC_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHIC_OM_V_readaddr,
        doutb     => AS_L2PHIC_OM_V_dout,
        sync_nent => AS_L2PHIC_OM_start,
        nent_o    => AS_L2PHIC_OM_AV_dout_nent
      );

    AS_L2PHIC_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHIC_OM_wea,
        addra     => AS_L2PHIC_OM_writeaddr,
        dina      => AS_L2PHIC_OM_din,
        wea_out       => AS_L2PHIC_OM_wea_delay,
        addra_out     => AS_L2PHIC_OM_writeaddr_delay,
        dina_out      => AS_L2PHIC_OM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHIC_OM_start
      );

    AS_L2PHID_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHID_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHID_BM_wea_delay,
        addra     => AS_L2PHID_BM_writeaddr_delay,
        dina      => AS_L2PHID_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHID_BM_V_readaddr,
        doutb     => AS_L2PHID_BM_V_dout,
        sync_nent => AS_L2PHID_BM_start,
        nent_o    => AS_L2PHID_BM_AV_dout_nent
      );

    AS_L2PHID_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHID_BM_wea,
        addra     => AS_L2PHID_BM_writeaddr,
        dina      => AS_L2PHID_BM_din,
        wea_out       => AS_L2PHID_BM_wea_delay,
        addra_out     => AS_L2PHID_BM_writeaddr_delay,
        dina_out      => AS_L2PHID_BM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHID_BM_start
      );

    AS_L2PHID_OM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L2PHID_OM"
      )
      port map (
        clka      => clk,
        wea       => AS_L2PHID_OM_wea_delay,
        addra     => AS_L2PHID_OM_writeaddr_delay,
        dina      => AS_L2PHID_OM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L2PHID_OM_V_readaddr,
        doutb     => AS_L2PHID_OM_V_dout,
        sync_nent => AS_L2PHID_OM_start,
        nent_o    => AS_L2PHID_OM_AV_dout_nent
      );

    AS_L2PHID_OM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L2PHID_OM_wea,
        addra     => AS_L2PHID_OM_writeaddr,
        dina      => AS_L2PHID_OM_din,
        wea_out       => AS_L2PHID_OM_wea_delay,
        addra_out     => AS_L2PHID_OM_writeaddr_delay,
        dina_out      => AS_L2PHID_OM_din_delay,
        done       => VMR_done,
        start      => AS_L2PHID_OM_start
      );

    AS_L3PHIA_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIA_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIA_BM_wea_delay,
        addra     => AS_L3PHIA_BM_writeaddr_delay,
        dina      => AS_L3PHIA_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIA_BM_V_readaddr,
        doutb     => AS_L3PHIA_BM_V_dout,
        sync_nent => AS_L3PHIA_BM_start,
        nent_o    => AS_L3PHIA_BM_AV_dout_nent
      );

    AS_L3PHIA_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIA_BM_wea,
        addra     => AS_L3PHIA_BM_writeaddr,
        dina      => AS_L3PHIA_BM_din,
        wea_out       => AS_L3PHIA_BM_wea_delay,
        addra_out     => AS_L3PHIA_BM_writeaddr_delay,
        dina_out      => AS_L3PHIA_BM_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIA_BM_start
      );

    AS_L3PHIB_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIB_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIB_BM_wea_delay,
        addra     => AS_L3PHIB_BM_writeaddr_delay,
        dina      => AS_L3PHIB_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIB_BM_V_readaddr,
        doutb     => AS_L3PHIB_BM_V_dout,
        sync_nent => AS_L3PHIB_BM_start,
        nent_o    => AS_L3PHIB_BM_AV_dout_nent
      );

    AS_L3PHIB_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIB_BM_wea,
        addra     => AS_L3PHIB_BM_writeaddr,
        dina      => AS_L3PHIB_BM_din,
        wea_out       => AS_L3PHIB_BM_wea_delay,
        addra_out     => AS_L3PHIB_BM_writeaddr_delay,
        dina_out      => AS_L3PHIB_BM_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIB_BM_start
      );

    AS_L3PHIB_BR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIB_BR"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIB_BR_wea_delay,
        addra     => AS_L3PHIB_BR_writeaddr_delay,
        dina      => AS_L3PHIB_BR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIB_BR_V_readaddr,
        doutb     => AS_L3PHIB_BR_V_dout,
        sync_nent => AS_L3PHIB_BR_start,
        nent_o    => AS_L3PHIB_BR_AV_dout_nent
      );

    AS_L3PHIB_BR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIB_BR_wea,
        addra     => AS_L3PHIB_BR_writeaddr,
        dina      => AS_L3PHIB_BR_din,
        wea_out       => AS_L3PHIB_BR_wea_delay,
        addra_out     => AS_L3PHIB_BR_writeaddr_delay,
        dina_out      => AS_L3PHIB_BR_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIB_BR_start
      );

    AS_L3PHIC_BL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIC_BL"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIC_BL_wea_delay,
        addra     => AS_L3PHIC_BL_writeaddr_delay,
        dina      => AS_L3PHIC_BL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIC_BL_V_readaddr,
        doutb     => AS_L3PHIC_BL_V_dout,
        sync_nent => AS_L3PHIC_BL_start,
        nent_o    => AS_L3PHIC_BL_AV_dout_nent
      );

    AS_L3PHIC_BL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIC_BL_wea,
        addra     => AS_L3PHIC_BL_writeaddr,
        dina      => AS_L3PHIC_BL_din,
        wea_out       => AS_L3PHIC_BL_wea_delay,
        addra_out     => AS_L3PHIC_BL_writeaddr_delay,
        dina_out      => AS_L3PHIC_BL_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIC_BL_start
      );

    AS_L3PHIC_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHIC_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHIC_BM_wea_delay,
        addra     => AS_L3PHIC_BM_writeaddr_delay,
        dina      => AS_L3PHIC_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHIC_BM_V_readaddr,
        doutb     => AS_L3PHIC_BM_V_dout,
        sync_nent => AS_L3PHIC_BM_start,
        nent_o    => AS_L3PHIC_BM_AV_dout_nent
      );

    AS_L3PHIC_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHIC_BM_wea,
        addra     => AS_L3PHIC_BM_writeaddr,
        dina      => AS_L3PHIC_BM_din,
        wea_out       => AS_L3PHIC_BM_wea_delay,
        addra_out     => AS_L3PHIC_BM_writeaddr_delay,
        dina_out      => AS_L3PHIC_BM_din_delay,
        done       => VMR_done,
        start      => AS_L3PHIC_BM_start
      );

    AS_L3PHID_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L3PHID_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L3PHID_BM_wea_delay,
        addra     => AS_L3PHID_BM_writeaddr_delay,
        dina      => AS_L3PHID_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L3PHID_BM_V_readaddr,
        doutb     => AS_L3PHID_BM_V_dout,
        sync_nent => AS_L3PHID_BM_start,
        nent_o    => AS_L3PHID_BM_AV_dout_nent
      );

    AS_L3PHID_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L3PHID_BM_wea,
        addra     => AS_L3PHID_BM_writeaddr,
        dina      => AS_L3PHID_BM_din,
        wea_out       => AS_L3PHID_BM_wea_delay,
        addra_out     => AS_L3PHID_BM_writeaddr_delay,
        dina_out      => AS_L3PHID_BM_din_delay,
        done       => VMR_done,
        start      => AS_L3PHID_BM_start
      );

    AS_L5PHIA_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIA_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIA_BM_wea_delay,
        addra     => AS_L5PHIA_BM_writeaddr_delay,
        dina      => AS_L5PHIA_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIA_BM_V_readaddr,
        doutb     => AS_L5PHIA_BM_V_dout,
        sync_nent => AS_L5PHIA_BM_start,
        nent_o    => AS_L5PHIA_BM_AV_dout_nent
      );

    AS_L5PHIA_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIA_BM_wea,
        addra     => AS_L5PHIA_BM_writeaddr,
        dina      => AS_L5PHIA_BM_din,
        wea_out       => AS_L5PHIA_BM_wea_delay,
        addra_out     => AS_L5PHIA_BM_writeaddr_delay,
        dina_out      => AS_L5PHIA_BM_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIA_BM_start
      );

    AS_L5PHIB_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIB_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIB_BM_wea_delay,
        addra     => AS_L5PHIB_BM_writeaddr_delay,
        dina      => AS_L5PHIB_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIB_BM_V_readaddr,
        doutb     => AS_L5PHIB_BM_V_dout,
        sync_nent => AS_L5PHIB_BM_start,
        nent_o    => AS_L5PHIB_BM_AV_dout_nent
      );

    AS_L5PHIB_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIB_BM_wea,
        addra     => AS_L5PHIB_BM_writeaddr,
        dina      => AS_L5PHIB_BM_din,
        wea_out       => AS_L5PHIB_BM_wea_delay,
        addra_out     => AS_L5PHIB_BM_writeaddr_delay,
        dina_out      => AS_L5PHIB_BM_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIB_BM_start
      );

    AS_L5PHIB_BR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIB_BR"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIB_BR_wea_delay,
        addra     => AS_L5PHIB_BR_writeaddr_delay,
        dina      => AS_L5PHIB_BR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIB_BR_V_readaddr,
        doutb     => AS_L5PHIB_BR_V_dout,
        sync_nent => AS_L5PHIB_BR_start,
        nent_o    => AS_L5PHIB_BR_AV_dout_nent
      );

    AS_L5PHIB_BR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIB_BR_wea,
        addra     => AS_L5PHIB_BR_writeaddr,
        dina      => AS_L5PHIB_BR_din,
        wea_out       => AS_L5PHIB_BR_wea_delay,
        addra_out     => AS_L5PHIB_BR_writeaddr_delay,
        dina_out      => AS_L5PHIB_BR_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIB_BR_start
      );

    AS_L5PHIC_BL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIC_BL"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIC_BL_wea_delay,
        addra     => AS_L5PHIC_BL_writeaddr_delay,
        dina      => AS_L5PHIC_BL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIC_BL_V_readaddr,
        doutb     => AS_L5PHIC_BL_V_dout,
        sync_nent => AS_L5PHIC_BL_start,
        nent_o    => AS_L5PHIC_BL_AV_dout_nent
      );

    AS_L5PHIC_BL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIC_BL_wea,
        addra     => AS_L5PHIC_BL_writeaddr,
        dina      => AS_L5PHIC_BL_din,
        wea_out       => AS_L5PHIC_BL_wea_delay,
        addra_out     => AS_L5PHIC_BL_writeaddr_delay,
        dina_out      => AS_L5PHIC_BL_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIC_BL_start
      );

    AS_L5PHIC_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHIC_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHIC_BM_wea_delay,
        addra     => AS_L5PHIC_BM_writeaddr_delay,
        dina      => AS_L5PHIC_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHIC_BM_V_readaddr,
        doutb     => AS_L5PHIC_BM_V_dout,
        sync_nent => AS_L5PHIC_BM_start,
        nent_o    => AS_L5PHIC_BM_AV_dout_nent
      );

    AS_L5PHIC_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHIC_BM_wea,
        addra     => AS_L5PHIC_BM_writeaddr,
        dina      => AS_L5PHIC_BM_din,
        wea_out       => AS_L5PHIC_BM_wea_delay,
        addra_out     => AS_L5PHIC_BM_writeaddr_delay,
        dina_out      => AS_L5PHIC_BM_din_delay,
        done       => VMR_done,
        start      => AS_L5PHIC_BM_start
      );

    AS_L5PHID_BM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_L5PHID_BM"
      )
      port map (
        clka      => clk,
        wea       => AS_L5PHID_BM_wea_delay,
        addra     => AS_L5PHID_BM_writeaddr_delay,
        dina      => AS_L5PHID_BM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_L5PHID_BM_V_readaddr,
        doutb     => AS_L5PHID_BM_V_dout,
        sync_nent => AS_L5PHID_BM_start,
        nent_o    => AS_L5PHID_BM_AV_dout_nent
      );

    AS_L5PHID_BM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_L5PHID_BM_wea,
        addra     => AS_L5PHID_BM_writeaddr,
        dina      => AS_L5PHID_BM_din,
        wea_out       => AS_L5PHID_BM_wea_delay,
        addra_out     => AS_L5PHID_BM_writeaddr_delay,
        dina_out      => AS_L5PHID_BM_din_delay,
        done       => VMR_done,
        start      => AS_L5PHID_BM_start
      );

    AS_D1PHIA_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIA_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIA_DM_wea_delay,
        addra     => AS_D1PHIA_DM_writeaddr_delay,
        dina      => AS_D1PHIA_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIA_DM_V_readaddr,
        doutb     => AS_D1PHIA_DM_V_dout,
        sync_nent => AS_D1PHIA_DM_start,
        nent_o    => AS_D1PHIA_DM_AV_dout_nent
      );

    AS_D1PHIA_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIA_DM_wea,
        addra     => AS_D1PHIA_DM_writeaddr,
        dina      => AS_D1PHIA_DM_din,
        wea_out       => AS_D1PHIA_DM_wea_delay,
        addra_out     => AS_D1PHIA_DM_writeaddr_delay,
        dina_out      => AS_D1PHIA_DM_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIA_DM_start
      );

    AS_D1PHIB_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIB_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIB_DM_wea_delay,
        addra     => AS_D1PHIB_DM_writeaddr_delay,
        dina      => AS_D1PHIB_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIB_DM_V_readaddr,
        doutb     => AS_D1PHIB_DM_V_dout,
        sync_nent => AS_D1PHIB_DM_start,
        nent_o    => AS_D1PHIB_DM_AV_dout_nent
      );

    AS_D1PHIB_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIB_DM_wea,
        addra     => AS_D1PHIB_DM_writeaddr,
        dina      => AS_D1PHIB_DM_din,
        wea_out       => AS_D1PHIB_DM_wea_delay,
        addra_out     => AS_D1PHIB_DM_writeaddr_delay,
        dina_out      => AS_D1PHIB_DM_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIB_DM_start
      );

    AS_D1PHIB_DR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIB_DR"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIB_DR_wea_delay,
        addra     => AS_D1PHIB_DR_writeaddr_delay,
        dina      => AS_D1PHIB_DR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIB_DR_V_readaddr,
        doutb     => AS_D1PHIB_DR_V_dout,
        sync_nent => AS_D1PHIB_DR_start,
        nent_o    => AS_D1PHIB_DR_AV_dout_nent
      );

    AS_D1PHIB_DR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIB_DR_wea,
        addra     => AS_D1PHIB_DR_writeaddr,
        dina      => AS_D1PHIB_DR_din,
        wea_out       => AS_D1PHIB_DR_wea_delay,
        addra_out     => AS_D1PHIB_DR_writeaddr_delay,
        dina_out      => AS_D1PHIB_DR_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIB_DR_start
      );

    AS_D1PHIC_DL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIC_DL"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIC_DL_wea_delay,
        addra     => AS_D1PHIC_DL_writeaddr_delay,
        dina      => AS_D1PHIC_DL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIC_DL_V_readaddr,
        doutb     => AS_D1PHIC_DL_V_dout,
        sync_nent => AS_D1PHIC_DL_start,
        nent_o    => AS_D1PHIC_DL_AV_dout_nent
      );

    AS_D1PHIC_DL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIC_DL_wea,
        addra     => AS_D1PHIC_DL_writeaddr,
        dina      => AS_D1PHIC_DL_din,
        wea_out       => AS_D1PHIC_DL_wea_delay,
        addra_out     => AS_D1PHIC_DL_writeaddr_delay,
        dina_out      => AS_D1PHIC_DL_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIC_DL_start
      );

    AS_D1PHIC_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHIC_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHIC_DM_wea_delay,
        addra     => AS_D1PHIC_DM_writeaddr_delay,
        dina      => AS_D1PHIC_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHIC_DM_V_readaddr,
        doutb     => AS_D1PHIC_DM_V_dout,
        sync_nent => AS_D1PHIC_DM_start,
        nent_o    => AS_D1PHIC_DM_AV_dout_nent
      );

    AS_D1PHIC_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHIC_DM_wea,
        addra     => AS_D1PHIC_DM_writeaddr,
        dina      => AS_D1PHIC_DM_din,
        wea_out       => AS_D1PHIC_DM_wea_delay,
        addra_out     => AS_D1PHIC_DM_writeaddr_delay,
        dina_out      => AS_D1PHIC_DM_din_delay,
        done       => VMR_done,
        start      => AS_D1PHIC_DM_start
      );

    AS_D1PHID_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D1PHID_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D1PHID_DM_wea_delay,
        addra     => AS_D1PHID_DM_writeaddr_delay,
        dina      => AS_D1PHID_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D1PHID_DM_V_readaddr,
        doutb     => AS_D1PHID_DM_V_dout,
        sync_nent => AS_D1PHID_DM_start,
        nent_o    => AS_D1PHID_DM_AV_dout_nent
      );

    AS_D1PHID_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D1PHID_DM_wea,
        addra     => AS_D1PHID_DM_writeaddr,
        dina      => AS_D1PHID_DM_din,
        wea_out       => AS_D1PHID_DM_wea_delay,
        addra_out     => AS_D1PHID_DM_writeaddr_delay,
        dina_out      => AS_D1PHID_DM_din_delay,
        done       => VMR_done,
        start      => AS_D1PHID_DM_start
      );

    AS_D3PHIA_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIA_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIA_DM_wea_delay,
        addra     => AS_D3PHIA_DM_writeaddr_delay,
        dina      => AS_D3PHIA_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIA_DM_V_readaddr,
        doutb     => AS_D3PHIA_DM_V_dout,
        sync_nent => AS_D3PHIA_DM_start,
        nent_o    => AS_D3PHIA_DM_AV_dout_nent
      );

    AS_D3PHIA_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIA_DM_wea,
        addra     => AS_D3PHIA_DM_writeaddr,
        dina      => AS_D3PHIA_DM_din,
        wea_out       => AS_D3PHIA_DM_wea_delay,
        addra_out     => AS_D3PHIA_DM_writeaddr_delay,
        dina_out      => AS_D3PHIA_DM_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIA_DM_start
      );

    AS_D3PHIB_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIB_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIB_DM_wea_delay,
        addra     => AS_D3PHIB_DM_writeaddr_delay,
        dina      => AS_D3PHIB_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIB_DM_V_readaddr,
        doutb     => AS_D3PHIB_DM_V_dout,
        sync_nent => AS_D3PHIB_DM_start,
        nent_o    => AS_D3PHIB_DM_AV_dout_nent
      );

    AS_D3PHIB_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIB_DM_wea,
        addra     => AS_D3PHIB_DM_writeaddr,
        dina      => AS_D3PHIB_DM_din,
        wea_out       => AS_D3PHIB_DM_wea_delay,
        addra_out     => AS_D3PHIB_DM_writeaddr_delay,
        dina_out      => AS_D3PHIB_DM_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIB_DM_start
      );

    AS_D3PHIB_DR : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIB_DR"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIB_DR_wea_delay,
        addra     => AS_D3PHIB_DR_writeaddr_delay,
        dina      => AS_D3PHIB_DR_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIB_DR_V_readaddr,
        doutb     => AS_D3PHIB_DR_V_dout,
        sync_nent => AS_D3PHIB_DR_start,
        nent_o    => AS_D3PHIB_DR_AV_dout_nent
      );

    AS_D3PHIB_DR_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIB_DR_wea,
        addra     => AS_D3PHIB_DR_writeaddr,
        dina      => AS_D3PHIB_DR_din,
        wea_out       => AS_D3PHIB_DR_wea_delay,
        addra_out     => AS_D3PHIB_DR_writeaddr_delay,
        dina_out      => AS_D3PHIB_DR_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIB_DR_start
      );

    AS_D3PHIC_DL : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIC_DL"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIC_DL_wea_delay,
        addra     => AS_D3PHIC_DL_writeaddr_delay,
        dina      => AS_D3PHIC_DL_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIC_DL_V_readaddr,
        doutb     => AS_D3PHIC_DL_V_dout,
        sync_nent => AS_D3PHIC_DL_start,
        nent_o    => AS_D3PHIC_DL_AV_dout_nent
      );

    AS_D3PHIC_DL_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIC_DL_wea,
        addra     => AS_D3PHIC_DL_writeaddr,
        dina      => AS_D3PHIC_DL_din,
        wea_out       => AS_D3PHIC_DL_wea_delay,
        addra_out     => AS_D3PHIC_DL_writeaddr_delay,
        dina_out      => AS_D3PHIC_DL_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIC_DL_start
      );

    AS_D3PHIC_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHIC_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHIC_DM_wea_delay,
        addra     => AS_D3PHIC_DM_writeaddr_delay,
        dina      => AS_D3PHIC_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHIC_DM_V_readaddr,
        doutb     => AS_D3PHIC_DM_V_dout,
        sync_nent => AS_D3PHIC_DM_start,
        nent_o    => AS_D3PHIC_DM_AV_dout_nent
      );

    AS_D3PHIC_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHIC_DM_wea,
        addra     => AS_D3PHIC_DM_writeaddr,
        dina      => AS_D3PHIC_DM_din,
        wea_out       => AS_D3PHIC_DM_wea_delay,
        addra_out     => AS_D3PHIC_DM_writeaddr_delay,
        dina_out      => AS_D3PHIC_DM_din_delay,
        done       => VMR_done,
        start      => AS_D3PHIC_DM_start
      );

    AS_D3PHID_DM : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 51,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "AS_D3PHID_DM"
      )
      port map (
        clka      => clk,
        wea       => AS_D3PHID_DM_wea_delay,
        addra     => AS_D3PHID_DM_writeaddr_delay,
        dina      => AS_D3PHID_DM_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => AS_D3PHID_DM_V_readaddr,
        doutb     => AS_D3PHID_DM_V_dout,
        sync_nent => AS_D3PHID_DM_start,
        nent_o    => AS_D3PHID_DM_AV_dout_nent
      );

    AS_D3PHID_DM_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_WIDTH       => 51
      )
      port map (
        clk      => clk,
        wea       => AS_D3PHID_DM_wea,
        addra     => AS_D3PHID_DM_writeaddr,
        dina      => AS_D3PHID_DM_din,
        wea_out       => AS_D3PHID_DM_wea_delay,
        addra_out     => AS_D3PHID_DM_writeaddr_delay,
        dina_out      => AS_D3PHID_DM_din_delay,
        done       => VMR_done,
        start      => AS_D3PHID_DM_start
      );

    VMSTE_L2PHIAn1_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIAn1_V_datatmp,
        dataout0 => VMSTE_L2PHIAn1_AV_dout(0),
        dataout1 => VMSTE_L2PHIAn1_AV_dout(1),
        dataout2 => VMSTE_L2PHIAn1_AV_dout(2),
        dataout3 => VMSTE_L2PHIAn1_AV_dout(3),
        dataout4 => VMSTE_L2PHIAn1_AV_dout(4)
      );

    VMSTE_L2PHIAn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIAn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIAn1_wea_delay,
        addra     => VMSTE_L2PHIAn1_writeaddr_delay,
        dina      => VMSTE_L2PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIAn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIAn1_AV_readaddr(4),VMSTE_L2PHIAn1_AV_readaddr(3),VMSTE_L2PHIAn1_AV_readaddr(2),VMSTE_L2PHIAn1_AV_readaddr(1),VMSTE_L2PHIAn1_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIAn1_V_datatmp,
        enb_nent  => VMSTE_L2PHIAn1_enb_nent,
        addr_nent  => VMSTE_L2PHIAn1_V_addr_nent,
        dout_nent  => VMSTE_L2PHIAn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIAn1_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIAn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIAn1_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIAn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIAn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIAn1_V_binmaskb
      );

    VMSTE_L2PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIAn1_wea,
        addra     => VMSTE_L2PHIAn1_writeaddr,
        dina      => VMSTE_L2PHIAn1_din,
        wea_out       => VMSTE_L2PHIAn1_wea_delay,
        addra_out     => VMSTE_L2PHIAn1_writeaddr_delay,
        dina_out      => VMSTE_L2PHIAn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIAn1_start
      );

    VMSTE_L2PHIAn2_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIAn2_V_datatmp,
        dataout0 => VMSTE_L2PHIAn2_AV_dout(0),
        dataout1 => VMSTE_L2PHIAn2_AV_dout(1),
        dataout2 => VMSTE_L2PHIAn2_AV_dout(2),
        dataout3 => VMSTE_L2PHIAn2_AV_dout(3),
        dataout4 => VMSTE_L2PHIAn2_AV_dout(4)
      );

    VMSTE_L2PHIAn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIAn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIAn2_wea_delay,
        addra     => VMSTE_L2PHIAn2_writeaddr_delay,
        dina      => VMSTE_L2PHIAn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIAn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIAn2_AV_readaddr(4),VMSTE_L2PHIAn2_AV_readaddr(3),VMSTE_L2PHIAn2_AV_readaddr(2),VMSTE_L2PHIAn2_AV_readaddr(1),VMSTE_L2PHIAn2_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIAn2_V_datatmp,
        enb_nent  => VMSTE_L2PHIAn2_enb_nent,
        addr_nent  => VMSTE_L2PHIAn2_V_addr_nent,
        dout_nent  => VMSTE_L2PHIAn2_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIAn2_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIAn2_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIAn2_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIAn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIAn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIAn2_V_binmaskb
      );

    VMSTE_L2PHIAn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIAn2_wea,
        addra     => VMSTE_L2PHIAn2_writeaddr,
        dina      => VMSTE_L2PHIAn2_din,
        wea_out       => VMSTE_L2PHIAn2_wea_delay,
        addra_out     => VMSTE_L2PHIAn2_writeaddr_delay,
        dina_out      => VMSTE_L2PHIAn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIAn2_start
      );

    VMSTE_L2PHIAn3_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIAn3_V_datatmp,
        dataout0 => VMSTE_L2PHIAn3_AV_dout(0),
        dataout1 => VMSTE_L2PHIAn3_AV_dout(1),
        dataout2 => VMSTE_L2PHIAn3_AV_dout(2),
        dataout3 => VMSTE_L2PHIAn3_AV_dout(3),
        dataout4 => VMSTE_L2PHIAn3_AV_dout(4)
      );

    VMSTE_L2PHIAn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIAn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIAn3_wea_delay,
        addra     => VMSTE_L2PHIAn3_writeaddr_delay,
        dina      => VMSTE_L2PHIAn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIAn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIAn3_AV_readaddr(4),VMSTE_L2PHIAn3_AV_readaddr(3),VMSTE_L2PHIAn3_AV_readaddr(2),VMSTE_L2PHIAn3_AV_readaddr(1),VMSTE_L2PHIAn3_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIAn3_V_datatmp,
        enb_nent  => VMSTE_L2PHIAn3_enb_nent,
        addr_nent  => VMSTE_L2PHIAn3_V_addr_nent,
        dout_nent  => VMSTE_L2PHIAn3_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIAn3_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIAn3_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIAn3_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIAn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIAn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIAn3_V_binmaskb
      );

    VMSTE_L2PHIAn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIAn3_wea,
        addra     => VMSTE_L2PHIAn3_writeaddr,
        dina      => VMSTE_L2PHIAn3_din,
        wea_out       => VMSTE_L2PHIAn3_wea_delay,
        addra_out     => VMSTE_L2PHIAn3_writeaddr_delay,
        dina_out      => VMSTE_L2PHIAn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIAn3_start
      );

    VMSTE_L2PHIBn1_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIBn1_V_datatmp,
        dataout0 => VMSTE_L2PHIBn1_AV_dout(0),
        dataout1 => VMSTE_L2PHIBn1_AV_dout(1),
        dataout2 => VMSTE_L2PHIBn1_AV_dout(2),
        dataout3 => VMSTE_L2PHIBn1_AV_dout(3),
        dataout4 => VMSTE_L2PHIBn1_AV_dout(4)
      );

    VMSTE_L2PHIBn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIBn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIBn1_wea_delay,
        addra     => VMSTE_L2PHIBn1_writeaddr_delay,
        dina      => VMSTE_L2PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIBn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIBn1_AV_readaddr(4),VMSTE_L2PHIBn1_AV_readaddr(3),VMSTE_L2PHIBn1_AV_readaddr(2),VMSTE_L2PHIBn1_AV_readaddr(1),VMSTE_L2PHIBn1_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIBn1_V_datatmp,
        enb_nent  => VMSTE_L2PHIBn1_enb_nent,
        addr_nent  => VMSTE_L2PHIBn1_V_addr_nent,
        dout_nent  => VMSTE_L2PHIBn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIBn1_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIBn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIBn1_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIBn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIBn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIBn1_V_binmaskb
      );

    VMSTE_L2PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIBn1_wea,
        addra     => VMSTE_L2PHIBn1_writeaddr,
        dina      => VMSTE_L2PHIBn1_din,
        wea_out       => VMSTE_L2PHIBn1_wea_delay,
        addra_out     => VMSTE_L2PHIBn1_writeaddr_delay,
        dina_out      => VMSTE_L2PHIBn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIBn1_start
      );

    VMSTE_L2PHIBn2_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIBn2_V_datatmp,
        dataout0 => VMSTE_L2PHIBn2_AV_dout(0),
        dataout1 => VMSTE_L2PHIBn2_AV_dout(1),
        dataout2 => VMSTE_L2PHIBn2_AV_dout(2),
        dataout3 => VMSTE_L2PHIBn2_AV_dout(3),
        dataout4 => VMSTE_L2PHIBn2_AV_dout(4)
      );

    VMSTE_L2PHIBn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIBn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIBn2_wea_delay,
        addra     => VMSTE_L2PHIBn2_writeaddr_delay,
        dina      => VMSTE_L2PHIBn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIBn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIBn2_AV_readaddr(4),VMSTE_L2PHIBn2_AV_readaddr(3),VMSTE_L2PHIBn2_AV_readaddr(2),VMSTE_L2PHIBn2_AV_readaddr(1),VMSTE_L2PHIBn2_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIBn2_V_datatmp,
        enb_nent  => VMSTE_L2PHIBn2_enb_nent,
        addr_nent  => VMSTE_L2PHIBn2_V_addr_nent,
        dout_nent  => VMSTE_L2PHIBn2_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIBn2_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIBn2_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIBn2_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIBn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIBn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIBn2_V_binmaskb
      );

    VMSTE_L2PHIBn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIBn2_wea,
        addra     => VMSTE_L2PHIBn2_writeaddr,
        dina      => VMSTE_L2PHIBn2_din,
        wea_out       => VMSTE_L2PHIBn2_wea_delay,
        addra_out     => VMSTE_L2PHIBn2_writeaddr_delay,
        dina_out      => VMSTE_L2PHIBn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIBn2_start
      );

    VMSTE_L2PHIBn3_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIBn3_V_datatmp,
        dataout0 => VMSTE_L2PHIBn3_AV_dout(0),
        dataout1 => VMSTE_L2PHIBn3_AV_dout(1),
        dataout2 => VMSTE_L2PHIBn3_AV_dout(2),
        dataout3 => VMSTE_L2PHIBn3_AV_dout(3),
        dataout4 => VMSTE_L2PHIBn3_AV_dout(4)
      );

    VMSTE_L2PHIBn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIBn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIBn3_wea_delay,
        addra     => VMSTE_L2PHIBn3_writeaddr_delay,
        dina      => VMSTE_L2PHIBn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIBn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIBn3_AV_readaddr(4),VMSTE_L2PHIBn3_AV_readaddr(3),VMSTE_L2PHIBn3_AV_readaddr(2),VMSTE_L2PHIBn3_AV_readaddr(1),VMSTE_L2PHIBn3_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIBn3_V_datatmp,
        enb_nent  => VMSTE_L2PHIBn3_enb_nent,
        addr_nent  => VMSTE_L2PHIBn3_V_addr_nent,
        dout_nent  => VMSTE_L2PHIBn3_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIBn3_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIBn3_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIBn3_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIBn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIBn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIBn3_V_binmaskb
      );

    VMSTE_L2PHIBn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIBn3_wea,
        addra     => VMSTE_L2PHIBn3_writeaddr,
        dina      => VMSTE_L2PHIBn3_din,
        wea_out       => VMSTE_L2PHIBn3_wea_delay,
        addra_out     => VMSTE_L2PHIBn3_writeaddr_delay,
        dina_out      => VMSTE_L2PHIBn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIBn3_start
      );

    VMSTE_L2PHICn1_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHICn1_V_datatmp,
        dataout0 => VMSTE_L2PHICn1_AV_dout(0),
        dataout1 => VMSTE_L2PHICn1_AV_dout(1),
        dataout2 => VMSTE_L2PHICn1_AV_dout(2),
        dataout3 => VMSTE_L2PHICn1_AV_dout(3),
        dataout4 => VMSTE_L2PHICn1_AV_dout(4)
      );

    VMSTE_L2PHICn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHICn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHICn1_wea_delay,
        addra     => VMSTE_L2PHICn1_writeaddr_delay,
        dina      => VMSTE_L2PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHICn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHICn1_AV_readaddr(4),VMSTE_L2PHICn1_AV_readaddr(3),VMSTE_L2PHICn1_AV_readaddr(2),VMSTE_L2PHICn1_AV_readaddr(1),VMSTE_L2PHICn1_AV_readaddr(0)),
        doutb     => VMSTE_L2PHICn1_V_datatmp,
        enb_nent  => VMSTE_L2PHICn1_enb_nent,
        addr_nent  => VMSTE_L2PHICn1_V_addr_nent,
        dout_nent  => VMSTE_L2PHICn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHICn1_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHICn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHICn1_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHICn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHICn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHICn1_V_binmaskb
      );

    VMSTE_L2PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHICn1_wea,
        addra     => VMSTE_L2PHICn1_writeaddr,
        dina      => VMSTE_L2PHICn1_din,
        wea_out       => VMSTE_L2PHICn1_wea_delay,
        addra_out     => VMSTE_L2PHICn1_writeaddr_delay,
        dina_out      => VMSTE_L2PHICn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHICn1_start
      );

    VMSTE_L2PHICn2_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHICn2_V_datatmp,
        dataout0 => VMSTE_L2PHICn2_AV_dout(0),
        dataout1 => VMSTE_L2PHICn2_AV_dout(1),
        dataout2 => VMSTE_L2PHICn2_AV_dout(2),
        dataout3 => VMSTE_L2PHICn2_AV_dout(3),
        dataout4 => VMSTE_L2PHICn2_AV_dout(4)
      );

    VMSTE_L2PHICn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHICn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHICn2_wea_delay,
        addra     => VMSTE_L2PHICn2_writeaddr_delay,
        dina      => VMSTE_L2PHICn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHICn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHICn2_AV_readaddr(4),VMSTE_L2PHICn2_AV_readaddr(3),VMSTE_L2PHICn2_AV_readaddr(2),VMSTE_L2PHICn2_AV_readaddr(1),VMSTE_L2PHICn2_AV_readaddr(0)),
        doutb     => VMSTE_L2PHICn2_V_datatmp,
        enb_nent  => VMSTE_L2PHICn2_enb_nent,
        addr_nent  => VMSTE_L2PHICn2_V_addr_nent,
        dout_nent  => VMSTE_L2PHICn2_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHICn2_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHICn2_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHICn2_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHICn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHICn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHICn2_V_binmaskb
      );

    VMSTE_L2PHICn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHICn2_wea,
        addra     => VMSTE_L2PHICn2_writeaddr,
        dina      => VMSTE_L2PHICn2_din,
        wea_out       => VMSTE_L2PHICn2_wea_delay,
        addra_out     => VMSTE_L2PHICn2_writeaddr_delay,
        dina_out      => VMSTE_L2PHICn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHICn2_start
      );

    VMSTE_L2PHICn3_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHICn3_V_datatmp,
        dataout0 => VMSTE_L2PHICn3_AV_dout(0),
        dataout1 => VMSTE_L2PHICn3_AV_dout(1),
        dataout2 => VMSTE_L2PHICn3_AV_dout(2),
        dataout3 => VMSTE_L2PHICn3_AV_dout(3),
        dataout4 => VMSTE_L2PHICn3_AV_dout(4)
      );

    VMSTE_L2PHICn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHICn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHICn3_wea_delay,
        addra     => VMSTE_L2PHICn3_writeaddr_delay,
        dina      => VMSTE_L2PHICn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHICn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHICn3_AV_readaddr(4),VMSTE_L2PHICn3_AV_readaddr(3),VMSTE_L2PHICn3_AV_readaddr(2),VMSTE_L2PHICn3_AV_readaddr(1),VMSTE_L2PHICn3_AV_readaddr(0)),
        doutb     => VMSTE_L2PHICn3_V_datatmp,
        enb_nent  => VMSTE_L2PHICn3_enb_nent,
        addr_nent  => VMSTE_L2PHICn3_V_addr_nent,
        dout_nent  => VMSTE_L2PHICn3_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHICn3_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHICn3_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHICn3_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHICn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHICn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHICn3_V_binmaskb
      );

    VMSTE_L2PHICn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHICn3_wea,
        addra     => VMSTE_L2PHICn3_writeaddr,
        dina      => VMSTE_L2PHICn3_din,
        wea_out       => VMSTE_L2PHICn3_wea_delay,
        addra_out     => VMSTE_L2PHICn3_writeaddr_delay,
        dina_out      => VMSTE_L2PHICn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHICn3_start
      );

    VMSTE_L2PHIDn1_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIDn1_V_datatmp,
        dataout0 => VMSTE_L2PHIDn1_AV_dout(0),
        dataout1 => VMSTE_L2PHIDn1_AV_dout(1),
        dataout2 => VMSTE_L2PHIDn1_AV_dout(2),
        dataout3 => VMSTE_L2PHIDn1_AV_dout(3),
        dataout4 => VMSTE_L2PHIDn1_AV_dout(4)
      );

    VMSTE_L2PHIDn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIDn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIDn1_wea_delay,
        addra     => VMSTE_L2PHIDn1_writeaddr_delay,
        dina      => VMSTE_L2PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIDn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIDn1_AV_readaddr(4),VMSTE_L2PHIDn1_AV_readaddr(3),VMSTE_L2PHIDn1_AV_readaddr(2),VMSTE_L2PHIDn1_AV_readaddr(1),VMSTE_L2PHIDn1_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIDn1_V_datatmp,
        enb_nent  => VMSTE_L2PHIDn1_enb_nent,
        addr_nent  => VMSTE_L2PHIDn1_V_addr_nent,
        dout_nent  => VMSTE_L2PHIDn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIDn1_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIDn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIDn1_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIDn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIDn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIDn1_V_binmaskb
      );

    VMSTE_L2PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIDn1_wea,
        addra     => VMSTE_L2PHIDn1_writeaddr,
        dina      => VMSTE_L2PHIDn1_din,
        wea_out       => VMSTE_L2PHIDn1_wea_delay,
        addra_out     => VMSTE_L2PHIDn1_writeaddr_delay,
        dina_out      => VMSTE_L2PHIDn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIDn1_start
      );

    VMSTE_L2PHIDn2_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIDn2_V_datatmp,
        dataout0 => VMSTE_L2PHIDn2_AV_dout(0),
        dataout1 => VMSTE_L2PHIDn2_AV_dout(1),
        dataout2 => VMSTE_L2PHIDn2_AV_dout(2),
        dataout3 => VMSTE_L2PHIDn2_AV_dout(3),
        dataout4 => VMSTE_L2PHIDn2_AV_dout(4)
      );

    VMSTE_L2PHIDn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIDn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIDn2_wea_delay,
        addra     => VMSTE_L2PHIDn2_writeaddr_delay,
        dina      => VMSTE_L2PHIDn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIDn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIDn2_AV_readaddr(4),VMSTE_L2PHIDn2_AV_readaddr(3),VMSTE_L2PHIDn2_AV_readaddr(2),VMSTE_L2PHIDn2_AV_readaddr(1),VMSTE_L2PHIDn2_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIDn2_V_datatmp,
        enb_nent  => VMSTE_L2PHIDn2_enb_nent,
        addr_nent  => VMSTE_L2PHIDn2_V_addr_nent,
        dout_nent  => VMSTE_L2PHIDn2_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIDn2_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIDn2_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIDn2_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIDn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIDn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIDn2_V_binmaskb
      );

    VMSTE_L2PHIDn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIDn2_wea,
        addra     => VMSTE_L2PHIDn2_writeaddr,
        dina      => VMSTE_L2PHIDn2_din,
        wea_out       => VMSTE_L2PHIDn2_wea_delay,
        addra_out     => VMSTE_L2PHIDn2_writeaddr_delay,
        dina_out      => VMSTE_L2PHIDn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIDn2_start
      );

    VMSTE_L2PHIDn3_dataformat : entity work.vmstub16dout5
      port map (
        datain => VMSTE_L2PHIDn3_V_datatmp,
        dataout0 => VMSTE_L2PHIDn3_AV_dout(0),
        dataout1 => VMSTE_L2PHIDn3_AV_dout(1),
        dataout2 => VMSTE_L2PHIDn3_AV_dout(2),
        dataout3 => VMSTE_L2PHIDn3_AV_dout(3),
        dataout4 => VMSTE_L2PHIDn3_AV_dout(4)
      );

    VMSTE_L2PHIDn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L2PHIDn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L2PHIDn3_wea_delay,
        addra     => VMSTE_L2PHIDn3_writeaddr_delay,
        dina      => VMSTE_L2PHIDn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L2PHIDn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L2PHIDn3_AV_readaddr(4),VMSTE_L2PHIDn3_AV_readaddr(3),VMSTE_L2PHIDn3_AV_readaddr(2),VMSTE_L2PHIDn3_AV_readaddr(1),VMSTE_L2PHIDn3_AV_readaddr(0)),
        doutb     => VMSTE_L2PHIDn3_V_datatmp,
        enb_nent  => VMSTE_L2PHIDn3_enb_nent,
        addr_nent  => VMSTE_L2PHIDn3_V_addr_nent,
        dout_nent  => VMSTE_L2PHIDn3_AV_dout_nent,
        enb_binmaska  => VMSTE_L2PHIDn3_enb_binmaska,
        addr_binmaska  => VMSTE_L2PHIDn3_V_addr_binmaska,
        binmaska_o  => VMSTE_L2PHIDn3_V_binmaska,
        enb_binmaskb  => VMSTE_L2PHIDn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_L2PHIDn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L2PHIDn3_V_binmaskb
      );

    VMSTE_L2PHIDn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L2PHIDn3_wea,
        addra     => VMSTE_L2PHIDn3_writeaddr,
        dina      => VMSTE_L2PHIDn3_din,
        wea_out       => VMSTE_L2PHIDn3_wea_delay,
        addra_out     => VMSTE_L2PHIDn3_writeaddr_delay,
        dina_out      => VMSTE_L2PHIDn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_L2PHIDn3_start
      );

    VMSTE_L3PHIIn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_L3PHIIn1_V_datatmp,
        dataout0 => VMSTE_L3PHIIn1_AV_dout(0),
        dataout1 => VMSTE_L3PHIIn1_AV_dout(1)
      );

    VMSTE_L3PHIIn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L3PHIIn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L3PHIIn1_wea_delay,
        addra     => VMSTE_L3PHIIn1_writeaddr_delay,
        dina      => VMSTE_L3PHIIn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L3PHIIn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L3PHIIn1_AV_readaddr(1),VMSTE_L3PHIIn1_AV_readaddr(0)),
        doutb     => VMSTE_L3PHIIn1_V_datatmp,
        enb_nent  => VMSTE_L3PHIIn1_enb_nent,
        addr_nent  => VMSTE_L3PHIIn1_V_addr_nent,
        dout_nent  => VMSTE_L3PHIIn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L3PHIIn1_enb_binmaska,
        addr_binmaska  => VMSTE_L3PHIIn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L3PHIIn1_V_binmaska,
        enb_binmaskb  => VMSTE_L3PHIIn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L3PHIIn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L3PHIIn1_V_binmaskb
      );

    VMSTE_L3PHIIn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L3PHIIn1_wea,
        addra     => VMSTE_L3PHIIn1_writeaddr,
        dina      => VMSTE_L3PHIIn1_din,
        wea_out       => VMSTE_L3PHIIn1_wea_delay,
        addra_out     => VMSTE_L3PHIIn1_writeaddr_delay,
        dina_out      => VMSTE_L3PHIIn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L3PHIIn1_start
      );

    VMSTE_L3PHIJn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_L3PHIJn1_V_datatmp,
        dataout0 => VMSTE_L3PHIJn1_AV_dout(0),
        dataout1 => VMSTE_L3PHIJn1_AV_dout(1)
      );

    VMSTE_L3PHIJn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L3PHIJn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L3PHIJn1_wea_delay,
        addra     => VMSTE_L3PHIJn1_writeaddr_delay,
        dina      => VMSTE_L3PHIJn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L3PHIJn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L3PHIJn1_AV_readaddr(1),VMSTE_L3PHIJn1_AV_readaddr(0)),
        doutb     => VMSTE_L3PHIJn1_V_datatmp,
        enb_nent  => VMSTE_L3PHIJn1_enb_nent,
        addr_nent  => VMSTE_L3PHIJn1_V_addr_nent,
        dout_nent  => VMSTE_L3PHIJn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L3PHIJn1_enb_binmaska,
        addr_binmaska  => VMSTE_L3PHIJn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L3PHIJn1_V_binmaska,
        enb_binmaskb  => VMSTE_L3PHIJn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L3PHIJn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L3PHIJn1_V_binmaskb
      );

    VMSTE_L3PHIJn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L3PHIJn1_wea,
        addra     => VMSTE_L3PHIJn1_writeaddr,
        dina      => VMSTE_L3PHIJn1_din,
        wea_out       => VMSTE_L3PHIJn1_wea_delay,
        addra_out     => VMSTE_L3PHIJn1_writeaddr_delay,
        dina_out      => VMSTE_L3PHIJn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L3PHIJn1_start
      );

    VMSTE_L3PHIKn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_L3PHIKn1_V_datatmp,
        dataout0 => VMSTE_L3PHIKn1_AV_dout(0),
        dataout1 => VMSTE_L3PHIKn1_AV_dout(1)
      );

    VMSTE_L3PHIKn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L3PHIKn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L3PHIKn1_wea_delay,
        addra     => VMSTE_L3PHIKn1_writeaddr_delay,
        dina      => VMSTE_L3PHIKn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L3PHIKn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L3PHIKn1_AV_readaddr(1),VMSTE_L3PHIKn1_AV_readaddr(0)),
        doutb     => VMSTE_L3PHIKn1_V_datatmp,
        enb_nent  => VMSTE_L3PHIKn1_enb_nent,
        addr_nent  => VMSTE_L3PHIKn1_V_addr_nent,
        dout_nent  => VMSTE_L3PHIKn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L3PHIKn1_enb_binmaska,
        addr_binmaska  => VMSTE_L3PHIKn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L3PHIKn1_V_binmaska,
        enb_binmaskb  => VMSTE_L3PHIKn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L3PHIKn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L3PHIKn1_V_binmaskb
      );

    VMSTE_L3PHIKn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L3PHIKn1_wea,
        addra     => VMSTE_L3PHIKn1_writeaddr,
        dina      => VMSTE_L3PHIKn1_din,
        wea_out       => VMSTE_L3PHIKn1_wea_delay,
        addra_out     => VMSTE_L3PHIKn1_writeaddr_delay,
        dina_out      => VMSTE_L3PHIKn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L3PHIKn1_start
      );

    VMSTE_L3PHILn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_L3PHILn1_V_datatmp,
        dataout0 => VMSTE_L3PHILn1_AV_dout(0),
        dataout1 => VMSTE_L3PHILn1_AV_dout(1)
      );

    VMSTE_L3PHILn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L3PHILn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L3PHILn1_wea_delay,
        addra     => VMSTE_L3PHILn1_writeaddr_delay,
        dina      => VMSTE_L3PHILn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L3PHILn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L3PHILn1_AV_readaddr(1),VMSTE_L3PHILn1_AV_readaddr(0)),
        doutb     => VMSTE_L3PHILn1_V_datatmp,
        enb_nent  => VMSTE_L3PHILn1_enb_nent,
        addr_nent  => VMSTE_L3PHILn1_V_addr_nent,
        dout_nent  => VMSTE_L3PHILn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L3PHILn1_enb_binmaska,
        addr_binmaska  => VMSTE_L3PHILn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L3PHILn1_V_binmaska,
        enb_binmaskb  => VMSTE_L3PHILn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L3PHILn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L3PHILn1_V_binmaskb
      );

    VMSTE_L3PHILn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L3PHILn1_wea,
        addra     => VMSTE_L3PHILn1_writeaddr,
        dina      => VMSTE_L3PHILn1_din,
        wea_out       => VMSTE_L3PHILn1_wea_delay,
        addra_out     => VMSTE_L3PHILn1_writeaddr_delay,
        dina_out      => VMSTE_L3PHILn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L3PHILn1_start
      );

    VMSTE_D2PHIAn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D2PHIAn1_V_datatmp,
        dataout0 => VMSTE_D2PHIAn1_AV_dout(0),
        dataout1 => VMSTE_D2PHIAn1_AV_dout(1),
        dataout2 => VMSTE_D2PHIAn1_AV_dout(2)
      );

    VMSTE_D2PHIAn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D2PHIAn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D2PHIAn1_wea_delay,
        addra     => VMSTE_D2PHIAn1_writeaddr_delay,
        dina      => VMSTE_D2PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D2PHIAn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D2PHIAn1_AV_readaddr(2),VMSTE_D2PHIAn1_AV_readaddr(1),VMSTE_D2PHIAn1_AV_readaddr(0)),
        doutb     => VMSTE_D2PHIAn1_V_datatmp,
        enb_nent  => VMSTE_D2PHIAn1_enb_nent,
        addr_nent  => VMSTE_D2PHIAn1_V_addr_nent,
        dout_nent  => VMSTE_D2PHIAn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D2PHIAn1_enb_binmaska,
        addr_binmaska  => VMSTE_D2PHIAn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D2PHIAn1_V_binmaska,
        enb_binmaskb  => VMSTE_D2PHIAn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D2PHIAn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D2PHIAn1_V_binmaskb
      );

    VMSTE_D2PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D2PHIAn1_wea,
        addra     => VMSTE_D2PHIAn1_writeaddr,
        dina      => VMSTE_D2PHIAn1_din,
        wea_out       => VMSTE_D2PHIAn1_wea_delay,
        addra_out     => VMSTE_D2PHIAn1_writeaddr_delay,
        dina_out      => VMSTE_D2PHIAn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D2PHIAn1_start
      );

    VMSTE_D2PHIBn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D2PHIBn1_V_datatmp,
        dataout0 => VMSTE_D2PHIBn1_AV_dout(0),
        dataout1 => VMSTE_D2PHIBn1_AV_dout(1),
        dataout2 => VMSTE_D2PHIBn1_AV_dout(2)
      );

    VMSTE_D2PHIBn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D2PHIBn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D2PHIBn1_wea_delay,
        addra     => VMSTE_D2PHIBn1_writeaddr_delay,
        dina      => VMSTE_D2PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D2PHIBn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D2PHIBn1_AV_readaddr(2),VMSTE_D2PHIBn1_AV_readaddr(1),VMSTE_D2PHIBn1_AV_readaddr(0)),
        doutb     => VMSTE_D2PHIBn1_V_datatmp,
        enb_nent  => VMSTE_D2PHIBn1_enb_nent,
        addr_nent  => VMSTE_D2PHIBn1_V_addr_nent,
        dout_nent  => VMSTE_D2PHIBn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D2PHIBn1_enb_binmaska,
        addr_binmaska  => VMSTE_D2PHIBn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D2PHIBn1_V_binmaska,
        enb_binmaskb  => VMSTE_D2PHIBn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D2PHIBn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D2PHIBn1_V_binmaskb
      );

    VMSTE_D2PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D2PHIBn1_wea,
        addra     => VMSTE_D2PHIBn1_writeaddr,
        dina      => VMSTE_D2PHIBn1_din,
        wea_out       => VMSTE_D2PHIBn1_wea_delay,
        addra_out     => VMSTE_D2PHIBn1_writeaddr_delay,
        dina_out      => VMSTE_D2PHIBn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D2PHIBn1_start
      );

    VMSTE_D2PHICn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D2PHICn1_V_datatmp,
        dataout0 => VMSTE_D2PHICn1_AV_dout(0),
        dataout1 => VMSTE_D2PHICn1_AV_dout(1),
        dataout2 => VMSTE_D2PHICn1_AV_dout(2)
      );

    VMSTE_D2PHICn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D2PHICn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D2PHICn1_wea_delay,
        addra     => VMSTE_D2PHICn1_writeaddr_delay,
        dina      => VMSTE_D2PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D2PHICn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D2PHICn1_AV_readaddr(2),VMSTE_D2PHICn1_AV_readaddr(1),VMSTE_D2PHICn1_AV_readaddr(0)),
        doutb     => VMSTE_D2PHICn1_V_datatmp,
        enb_nent  => VMSTE_D2PHICn1_enb_nent,
        addr_nent  => VMSTE_D2PHICn1_V_addr_nent,
        dout_nent  => VMSTE_D2PHICn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D2PHICn1_enb_binmaska,
        addr_binmaska  => VMSTE_D2PHICn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D2PHICn1_V_binmaska,
        enb_binmaskb  => VMSTE_D2PHICn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D2PHICn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D2PHICn1_V_binmaskb
      );

    VMSTE_D2PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D2PHICn1_wea,
        addra     => VMSTE_D2PHICn1_writeaddr,
        dina      => VMSTE_D2PHICn1_din,
        wea_out       => VMSTE_D2PHICn1_wea_delay,
        addra_out     => VMSTE_D2PHICn1_writeaddr_delay,
        dina_out      => VMSTE_D2PHICn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D2PHICn1_start
      );

    VMSTE_D2PHIDn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D2PHIDn1_V_datatmp,
        dataout0 => VMSTE_D2PHIDn1_AV_dout(0),
        dataout1 => VMSTE_D2PHIDn1_AV_dout(1),
        dataout2 => VMSTE_D2PHIDn1_AV_dout(2)
      );

    VMSTE_D2PHIDn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D2PHIDn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D2PHIDn1_wea_delay,
        addra     => VMSTE_D2PHIDn1_writeaddr_delay,
        dina      => VMSTE_D2PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D2PHIDn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D2PHIDn1_AV_readaddr(2),VMSTE_D2PHIDn1_AV_readaddr(1),VMSTE_D2PHIDn1_AV_readaddr(0)),
        doutb     => VMSTE_D2PHIDn1_V_datatmp,
        enb_nent  => VMSTE_D2PHIDn1_enb_nent,
        addr_nent  => VMSTE_D2PHIDn1_V_addr_nent,
        dout_nent  => VMSTE_D2PHIDn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D2PHIDn1_enb_binmaska,
        addr_binmaska  => VMSTE_D2PHIDn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D2PHIDn1_V_binmaska,
        enb_binmaskb  => VMSTE_D2PHIDn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D2PHIDn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D2PHIDn1_V_binmaskb
      );

    VMSTE_D2PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D2PHIDn1_wea,
        addra     => VMSTE_D2PHIDn1_writeaddr,
        dina      => VMSTE_D2PHIDn1_din,
        wea_out       => VMSTE_D2PHIDn1_wea_delay,
        addra_out     => VMSTE_D2PHIDn1_writeaddr_delay,
        dina_out      => VMSTE_D2PHIDn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D2PHIDn1_start
      );

    VMSTE_D4PHIAn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D4PHIAn1_V_datatmp,
        dataout0 => VMSTE_D4PHIAn1_AV_dout(0),
        dataout1 => VMSTE_D4PHIAn1_AV_dout(1)
      );

    VMSTE_D4PHIAn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D4PHIAn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D4PHIAn1_wea_delay,
        addra     => VMSTE_D4PHIAn1_writeaddr_delay,
        dina      => VMSTE_D4PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D4PHIAn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D4PHIAn1_AV_readaddr(1),VMSTE_D4PHIAn1_AV_readaddr(0)),
        doutb     => VMSTE_D4PHIAn1_V_datatmp,
        enb_nent  => VMSTE_D4PHIAn1_enb_nent,
        addr_nent  => VMSTE_D4PHIAn1_V_addr_nent,
        dout_nent  => VMSTE_D4PHIAn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D4PHIAn1_enb_binmaska,
        addr_binmaska  => VMSTE_D4PHIAn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D4PHIAn1_V_binmaska,
        enb_binmaskb  => VMSTE_D4PHIAn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D4PHIAn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D4PHIAn1_V_binmaskb
      );

    VMSTE_D4PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D4PHIAn1_wea,
        addra     => VMSTE_D4PHIAn1_writeaddr,
        dina      => VMSTE_D4PHIAn1_din,
        wea_out       => VMSTE_D4PHIAn1_wea_delay,
        addra_out     => VMSTE_D4PHIAn1_writeaddr_delay,
        dina_out      => VMSTE_D4PHIAn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D4PHIAn1_start
      );

    VMSTE_D4PHIBn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D4PHIBn1_V_datatmp,
        dataout0 => VMSTE_D4PHIBn1_AV_dout(0),
        dataout1 => VMSTE_D4PHIBn1_AV_dout(1)
      );

    VMSTE_D4PHIBn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D4PHIBn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D4PHIBn1_wea_delay,
        addra     => VMSTE_D4PHIBn1_writeaddr_delay,
        dina      => VMSTE_D4PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D4PHIBn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D4PHIBn1_AV_readaddr(1),VMSTE_D4PHIBn1_AV_readaddr(0)),
        doutb     => VMSTE_D4PHIBn1_V_datatmp,
        enb_nent  => VMSTE_D4PHIBn1_enb_nent,
        addr_nent  => VMSTE_D4PHIBn1_V_addr_nent,
        dout_nent  => VMSTE_D4PHIBn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D4PHIBn1_enb_binmaska,
        addr_binmaska  => VMSTE_D4PHIBn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D4PHIBn1_V_binmaska,
        enb_binmaskb  => VMSTE_D4PHIBn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D4PHIBn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D4PHIBn1_V_binmaskb
      );

    VMSTE_D4PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D4PHIBn1_wea,
        addra     => VMSTE_D4PHIBn1_writeaddr,
        dina      => VMSTE_D4PHIBn1_din,
        wea_out       => VMSTE_D4PHIBn1_wea_delay,
        addra_out     => VMSTE_D4PHIBn1_writeaddr_delay,
        dina_out      => VMSTE_D4PHIBn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D4PHIBn1_start
      );

    VMSTE_D4PHICn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D4PHICn1_V_datatmp,
        dataout0 => VMSTE_D4PHICn1_AV_dout(0),
        dataout1 => VMSTE_D4PHICn1_AV_dout(1)
      );

    VMSTE_D4PHICn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D4PHICn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D4PHICn1_wea_delay,
        addra     => VMSTE_D4PHICn1_writeaddr_delay,
        dina      => VMSTE_D4PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D4PHICn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D4PHICn1_AV_readaddr(1),VMSTE_D4PHICn1_AV_readaddr(0)),
        doutb     => VMSTE_D4PHICn1_V_datatmp,
        enb_nent  => VMSTE_D4PHICn1_enb_nent,
        addr_nent  => VMSTE_D4PHICn1_V_addr_nent,
        dout_nent  => VMSTE_D4PHICn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D4PHICn1_enb_binmaska,
        addr_binmaska  => VMSTE_D4PHICn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D4PHICn1_V_binmaska,
        enb_binmaskb  => VMSTE_D4PHICn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D4PHICn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D4PHICn1_V_binmaskb
      );

    VMSTE_D4PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D4PHICn1_wea,
        addra     => VMSTE_D4PHICn1_writeaddr,
        dina      => VMSTE_D4PHICn1_din,
        wea_out       => VMSTE_D4PHICn1_wea_delay,
        addra_out     => VMSTE_D4PHICn1_writeaddr_delay,
        dina_out      => VMSTE_D4PHICn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D4PHICn1_start
      );

    VMSTE_D4PHIDn1_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D4PHIDn1_V_datatmp,
        dataout0 => VMSTE_D4PHIDn1_AV_dout(0),
        dataout1 => VMSTE_D4PHIDn1_AV_dout(1)
      );

    VMSTE_D4PHIDn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D4PHIDn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D4PHIDn1_wea_delay,
        addra     => VMSTE_D4PHIDn1_writeaddr_delay,
        dina      => VMSTE_D4PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D4PHIDn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D4PHIDn1_AV_readaddr(1),VMSTE_D4PHIDn1_AV_readaddr(0)),
        doutb     => VMSTE_D4PHIDn1_V_datatmp,
        enb_nent  => VMSTE_D4PHIDn1_enb_nent,
        addr_nent  => VMSTE_D4PHIDn1_V_addr_nent,
        dout_nent  => VMSTE_D4PHIDn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D4PHIDn1_enb_binmaska,
        addr_binmaska  => VMSTE_D4PHIDn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D4PHIDn1_V_binmaska,
        enb_binmaskb  => VMSTE_D4PHIDn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D4PHIDn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D4PHIDn1_V_binmaskb
      );

    VMSTE_D4PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D4PHIDn1_wea,
        addra     => VMSTE_D4PHIDn1_writeaddr,
        dina      => VMSTE_D4PHIDn1_din,
        wea_out       => VMSTE_D4PHIDn1_wea_delay,
        addra_out     => VMSTE_D4PHIDn1_writeaddr_delay,
        dina_out      => VMSTE_D4PHIDn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D4PHIDn1_start
      );

    VMSTE_D1PHIXn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIXn1_V_datatmp,
        dataout0 => VMSTE_D1PHIXn1_AV_dout(0),
        dataout1 => VMSTE_D1PHIXn1_AV_dout(1),
        dataout2 => VMSTE_D1PHIXn1_AV_dout(2)
      );

    VMSTE_D1PHIXn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIXn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIXn1_wea_delay,
        addra     => VMSTE_D1PHIXn1_writeaddr_delay,
        dina      => VMSTE_D1PHIXn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIXn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIXn1_AV_readaddr(2),VMSTE_D1PHIXn1_AV_readaddr(1),VMSTE_D1PHIXn1_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIXn1_V_datatmp,
        enb_nent  => VMSTE_D1PHIXn1_enb_nent,
        addr_nent  => VMSTE_D1PHIXn1_V_addr_nent,
        dout_nent  => VMSTE_D1PHIXn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIXn1_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIXn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIXn1_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIXn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIXn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIXn1_V_binmaskb
      );

    VMSTE_D1PHIXn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIXn1_wea,
        addra     => VMSTE_D1PHIXn1_writeaddr,
        dina      => VMSTE_D1PHIXn1_din,
        wea_out       => VMSTE_D1PHIXn1_wea_delay,
        addra_out     => VMSTE_D1PHIXn1_writeaddr_delay,
        dina_out      => VMSTE_D1PHIXn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIXn1_start
      );

    VMSTE_D1PHIXn2_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIXn2_V_datatmp,
        dataout0 => VMSTE_D1PHIXn2_AV_dout(0),
        dataout1 => VMSTE_D1PHIXn2_AV_dout(1),
        dataout2 => VMSTE_D1PHIXn2_AV_dout(2)
      );

    VMSTE_D1PHIXn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIXn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIXn2_wea_delay,
        addra     => VMSTE_D1PHIXn2_writeaddr_delay,
        dina      => VMSTE_D1PHIXn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIXn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIXn2_AV_readaddr(2),VMSTE_D1PHIXn2_AV_readaddr(1),VMSTE_D1PHIXn2_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIXn2_V_datatmp,
        enb_nent  => VMSTE_D1PHIXn2_enb_nent,
        addr_nent  => VMSTE_D1PHIXn2_V_addr_nent,
        dout_nent  => VMSTE_D1PHIXn2_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIXn2_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIXn2_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIXn2_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIXn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIXn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIXn2_V_binmaskb
      );

    VMSTE_D1PHIXn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIXn2_wea,
        addra     => VMSTE_D1PHIXn2_writeaddr,
        dina      => VMSTE_D1PHIXn2_din,
        wea_out       => VMSTE_D1PHIXn2_wea_delay,
        addra_out     => VMSTE_D1PHIXn2_writeaddr_delay,
        dina_out      => VMSTE_D1PHIXn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIXn2_start
      );

    VMSTE_D1PHIYn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIYn1_V_datatmp,
        dataout0 => VMSTE_D1PHIYn1_AV_dout(0),
        dataout1 => VMSTE_D1PHIYn1_AV_dout(1),
        dataout2 => VMSTE_D1PHIYn1_AV_dout(2)
      );

    VMSTE_D1PHIYn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIYn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIYn1_wea_delay,
        addra     => VMSTE_D1PHIYn1_writeaddr_delay,
        dina      => VMSTE_D1PHIYn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIYn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIYn1_AV_readaddr(2),VMSTE_D1PHIYn1_AV_readaddr(1),VMSTE_D1PHIYn1_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIYn1_V_datatmp,
        enb_nent  => VMSTE_D1PHIYn1_enb_nent,
        addr_nent  => VMSTE_D1PHIYn1_V_addr_nent,
        dout_nent  => VMSTE_D1PHIYn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIYn1_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIYn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIYn1_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIYn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIYn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIYn1_V_binmaskb
      );

    VMSTE_D1PHIYn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIYn1_wea,
        addra     => VMSTE_D1PHIYn1_writeaddr,
        dina      => VMSTE_D1PHIYn1_din,
        wea_out       => VMSTE_D1PHIYn1_wea_delay,
        addra_out     => VMSTE_D1PHIYn1_writeaddr_delay,
        dina_out      => VMSTE_D1PHIYn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIYn1_start
      );

    VMSTE_D1PHIYn2_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIYn2_V_datatmp,
        dataout0 => VMSTE_D1PHIYn2_AV_dout(0),
        dataout1 => VMSTE_D1PHIYn2_AV_dout(1),
        dataout2 => VMSTE_D1PHIYn2_AV_dout(2)
      );

    VMSTE_D1PHIYn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIYn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIYn2_wea_delay,
        addra     => VMSTE_D1PHIYn2_writeaddr_delay,
        dina      => VMSTE_D1PHIYn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIYn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIYn2_AV_readaddr(2),VMSTE_D1PHIYn2_AV_readaddr(1),VMSTE_D1PHIYn2_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIYn2_V_datatmp,
        enb_nent  => VMSTE_D1PHIYn2_enb_nent,
        addr_nent  => VMSTE_D1PHIYn2_V_addr_nent,
        dout_nent  => VMSTE_D1PHIYn2_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIYn2_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIYn2_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIYn2_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIYn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIYn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIYn2_V_binmaskb
      );

    VMSTE_D1PHIYn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIYn2_wea,
        addra     => VMSTE_D1PHIYn2_writeaddr,
        dina      => VMSTE_D1PHIYn2_din,
        wea_out       => VMSTE_D1PHIYn2_wea_delay,
        addra_out     => VMSTE_D1PHIYn2_writeaddr_delay,
        dina_out      => VMSTE_D1PHIYn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIYn2_start
      );

    VMSTE_D1PHIZn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIZn1_V_datatmp,
        dataout0 => VMSTE_D1PHIZn1_AV_dout(0),
        dataout1 => VMSTE_D1PHIZn1_AV_dout(1),
        dataout2 => VMSTE_D1PHIZn1_AV_dout(2)
      );

    VMSTE_D1PHIZn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIZn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIZn1_wea_delay,
        addra     => VMSTE_D1PHIZn1_writeaddr_delay,
        dina      => VMSTE_D1PHIZn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIZn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIZn1_AV_readaddr(2),VMSTE_D1PHIZn1_AV_readaddr(1),VMSTE_D1PHIZn1_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIZn1_V_datatmp,
        enb_nent  => VMSTE_D1PHIZn1_enb_nent,
        addr_nent  => VMSTE_D1PHIZn1_V_addr_nent,
        dout_nent  => VMSTE_D1PHIZn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIZn1_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIZn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIZn1_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIZn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIZn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIZn1_V_binmaskb
      );

    VMSTE_D1PHIZn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIZn1_wea,
        addra     => VMSTE_D1PHIZn1_writeaddr,
        dina      => VMSTE_D1PHIZn1_din,
        wea_out       => VMSTE_D1PHIZn1_wea_delay,
        addra_out     => VMSTE_D1PHIZn1_writeaddr_delay,
        dina_out      => VMSTE_D1PHIZn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIZn1_start
      );

    VMSTE_D1PHIZn2_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIZn2_V_datatmp,
        dataout0 => VMSTE_D1PHIZn2_AV_dout(0),
        dataout1 => VMSTE_D1PHIZn2_AV_dout(1),
        dataout2 => VMSTE_D1PHIZn2_AV_dout(2)
      );

    VMSTE_D1PHIZn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIZn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIZn2_wea_delay,
        addra     => VMSTE_D1PHIZn2_writeaddr_delay,
        dina      => VMSTE_D1PHIZn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIZn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIZn2_AV_readaddr(2),VMSTE_D1PHIZn2_AV_readaddr(1),VMSTE_D1PHIZn2_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIZn2_V_datatmp,
        enb_nent  => VMSTE_D1PHIZn2_enb_nent,
        addr_nent  => VMSTE_D1PHIZn2_V_addr_nent,
        dout_nent  => VMSTE_D1PHIZn2_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIZn2_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIZn2_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIZn2_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIZn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIZn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIZn2_V_binmaskb
      );

    VMSTE_D1PHIZn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIZn2_wea,
        addra     => VMSTE_D1PHIZn2_writeaddr,
        dina      => VMSTE_D1PHIZn2_din,
        wea_out       => VMSTE_D1PHIZn2_wea_delay,
        addra_out     => VMSTE_D1PHIZn2_writeaddr_delay,
        dina_out      => VMSTE_D1PHIZn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIZn2_start
      );

    VMSTE_D1PHIWn1_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIWn1_V_datatmp,
        dataout0 => VMSTE_D1PHIWn1_AV_dout(0),
        dataout1 => VMSTE_D1PHIWn1_AV_dout(1),
        dataout2 => VMSTE_D1PHIWn1_AV_dout(2)
      );

    VMSTE_D1PHIWn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIWn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIWn1_wea_delay,
        addra     => VMSTE_D1PHIWn1_writeaddr_delay,
        dina      => VMSTE_D1PHIWn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIWn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIWn1_AV_readaddr(2),VMSTE_D1PHIWn1_AV_readaddr(1),VMSTE_D1PHIWn1_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIWn1_V_datatmp,
        enb_nent  => VMSTE_D1PHIWn1_enb_nent,
        addr_nent  => VMSTE_D1PHIWn1_V_addr_nent,
        dout_nent  => VMSTE_D1PHIWn1_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIWn1_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIWn1_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIWn1_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIWn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIWn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIWn1_V_binmaskb
      );

    VMSTE_D1PHIWn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIWn1_wea,
        addra     => VMSTE_D1PHIWn1_writeaddr,
        dina      => VMSTE_D1PHIWn1_din,
        wea_out       => VMSTE_D1PHIWn1_wea_delay,
        addra_out     => VMSTE_D1PHIWn1_writeaddr_delay,
        dina_out      => VMSTE_D1PHIWn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIWn1_start
      );

    VMSTE_D1PHIWn2_dataformat : entity work.vmstub16dout3
      port map (
        datain => VMSTE_D1PHIWn2_V_datatmp,
        dataout0 => VMSTE_D1PHIWn2_AV_dout(0),
        dataout1 => VMSTE_D1PHIWn2_AV_dout(1),
        dataout2 => VMSTE_D1PHIWn2_AV_dout(2)
      );

    VMSTE_D1PHIWn2 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIWn2",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIWn2_wea_delay,
        addra     => VMSTE_D1PHIWn2_writeaddr_delay,
        dina      => VMSTE_D1PHIWn2_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIWn2_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIWn2_AV_readaddr(2),VMSTE_D1PHIWn2_AV_readaddr(1),VMSTE_D1PHIWn2_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIWn2_V_datatmp,
        enb_nent  => VMSTE_D1PHIWn2_enb_nent,
        addr_nent  => VMSTE_D1PHIWn2_V_addr_nent,
        dout_nent  => VMSTE_D1PHIWn2_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIWn2_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIWn2_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIWn2_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIWn2_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIWn2_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIWn2_V_binmaskb
      );

    VMSTE_D1PHIWn2_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIWn2_wea,
        addra     => VMSTE_D1PHIWn2_writeaddr,
        dina      => VMSTE_D1PHIWn2_din,
        wea_out       => VMSTE_D1PHIWn2_wea_delay,
        addra_out     => VMSTE_D1PHIWn2_writeaddr_delay,
        dina_out      => VMSTE_D1PHIWn2_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIWn2_start
      );

    VMSTE_D1PHIXn3_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D1PHIXn3_V_datatmp,
        dataout0 => VMSTE_D1PHIXn3_AV_dout(0),
        dataout1 => VMSTE_D1PHIXn3_AV_dout(1)
      );

    VMSTE_D1PHIXn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIXn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIXn3_wea_delay,
        addra     => VMSTE_D1PHIXn3_writeaddr_delay,
        dina      => VMSTE_D1PHIXn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIXn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIXn3_AV_readaddr(1),VMSTE_D1PHIXn3_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIXn3_V_datatmp,
        enb_nent  => VMSTE_D1PHIXn3_enb_nent,
        addr_nent  => VMSTE_D1PHIXn3_V_addr_nent,
        dout_nent  => VMSTE_D1PHIXn3_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIXn3_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIXn3_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIXn3_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIXn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIXn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIXn3_V_binmaskb
      );

    VMSTE_D1PHIXn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIXn3_wea,
        addra     => VMSTE_D1PHIXn3_writeaddr,
        dina      => VMSTE_D1PHIXn3_din,
        wea_out       => VMSTE_D1PHIXn3_wea_delay,
        addra_out     => VMSTE_D1PHIXn3_writeaddr_delay,
        dina_out      => VMSTE_D1PHIXn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIXn3_start
      );

    VMSTE_D1PHIYn3_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D1PHIYn3_V_datatmp,
        dataout0 => VMSTE_D1PHIYn3_AV_dout(0),
        dataout1 => VMSTE_D1PHIYn3_AV_dout(1)
      );

    VMSTE_D1PHIYn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIYn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIYn3_wea_delay,
        addra     => VMSTE_D1PHIYn3_writeaddr_delay,
        dina      => VMSTE_D1PHIYn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIYn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIYn3_AV_readaddr(1),VMSTE_D1PHIYn3_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIYn3_V_datatmp,
        enb_nent  => VMSTE_D1PHIYn3_enb_nent,
        addr_nent  => VMSTE_D1PHIYn3_V_addr_nent,
        dout_nent  => VMSTE_D1PHIYn3_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIYn3_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIYn3_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIYn3_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIYn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIYn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIYn3_V_binmaskb
      );

    VMSTE_D1PHIYn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIYn3_wea,
        addra     => VMSTE_D1PHIYn3_writeaddr,
        dina      => VMSTE_D1PHIYn3_din,
        wea_out       => VMSTE_D1PHIYn3_wea_delay,
        addra_out     => VMSTE_D1PHIYn3_writeaddr_delay,
        dina_out      => VMSTE_D1PHIYn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIYn3_start
      );

    VMSTE_D1PHIZn3_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D1PHIZn3_V_datatmp,
        dataout0 => VMSTE_D1PHIZn3_AV_dout(0),
        dataout1 => VMSTE_D1PHIZn3_AV_dout(1)
      );

    VMSTE_D1PHIZn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIZn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIZn3_wea_delay,
        addra     => VMSTE_D1PHIZn3_writeaddr_delay,
        dina      => VMSTE_D1PHIZn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIZn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIZn3_AV_readaddr(1),VMSTE_D1PHIZn3_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIZn3_V_datatmp,
        enb_nent  => VMSTE_D1PHIZn3_enb_nent,
        addr_nent  => VMSTE_D1PHIZn3_V_addr_nent,
        dout_nent  => VMSTE_D1PHIZn3_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIZn3_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIZn3_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIZn3_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIZn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIZn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIZn3_V_binmaskb
      );

    VMSTE_D1PHIZn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIZn3_wea,
        addra     => VMSTE_D1PHIZn3_writeaddr,
        dina      => VMSTE_D1PHIZn3_din,
        wea_out       => VMSTE_D1PHIZn3_wea_delay,
        addra_out     => VMSTE_D1PHIZn3_writeaddr_delay,
        dina_out      => VMSTE_D1PHIZn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIZn3_start
      );

    VMSTE_D1PHIWn3_dataformat : entity work.vmstub16dout2
      port map (
        datain => VMSTE_D1PHIWn3_V_datatmp,
        dataout0 => VMSTE_D1PHIWn3_AV_dout(0),
        dataout1 => VMSTE_D1PHIWn3_AV_dout(1)
      );

    VMSTE_D1PHIWn3 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 16,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_D1PHIWn3",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 2
      )
      port map (
        clka      => clk,
        wea       => VMSTE_D1PHIWn3_wea_delay,
        addra     => VMSTE_D1PHIWn3_writeaddr_delay,
        dina      => VMSTE_D1PHIWn3_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_D1PHIWn3_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_D1PHIWn3_AV_readaddr(1),VMSTE_D1PHIWn3_AV_readaddr(0)),
        doutb     => VMSTE_D1PHIWn3_V_datatmp,
        enb_nent  => VMSTE_D1PHIWn3_enb_nent,
        addr_nent  => VMSTE_D1PHIWn3_V_addr_nent,
        dout_nent  => VMSTE_D1PHIWn3_AV_dout_nent,
        enb_binmaska  => VMSTE_D1PHIWn3_enb_binmaska,
        addr_binmaska  => VMSTE_D1PHIWn3_V_addr_binmaska,
        binmaska_o  => VMSTE_D1PHIWn3_V_binmaska,
        enb_binmaskb  => VMSTE_D1PHIWn3_enb_binmaskb,
        addr_binmaskb  => VMSTE_D1PHIWn3_V_addr_binmaskb,
        binmaskb_o  => VMSTE_D1PHIWn3_V_binmaskb
      );

    VMSTE_D1PHIWn3_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 16
      )
      port map (
        clk      => clk,
        wea       => VMSTE_D1PHIWn3_wea,
        addra     => VMSTE_D1PHIWn3_writeaddr,
        dina      => VMSTE_D1PHIWn3_din,
        wea_out       => VMSTE_D1PHIWn3_wea_delay,
        addra_out     => VMSTE_D1PHIWn3_writeaddr_delay,
        dina_out      => VMSTE_D1PHIWn3_din_delay,
        done       => VMR_done,
        start      => VMSTE_D1PHIWn3_start
      );

    VMSTE_L4PHIAn1_dataformat : entity work.vmstub17dout5
      port map (
        datain => VMSTE_L4PHIAn1_V_datatmp,
        dataout0 => VMSTE_L4PHIAn1_AV_dout(0),
        dataout1 => VMSTE_L4PHIAn1_AV_dout(1),
        dataout2 => VMSTE_L4PHIAn1_AV_dout(2),
        dataout3 => VMSTE_L4PHIAn1_AV_dout(3),
        dataout4 => VMSTE_L4PHIAn1_AV_dout(4)
      );

    VMSTE_L4PHIAn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L4PHIAn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L4PHIAn1_wea_delay,
        addra     => VMSTE_L4PHIAn1_writeaddr_delay,
        dina      => VMSTE_L4PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L4PHIAn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L4PHIAn1_AV_readaddr(4),VMSTE_L4PHIAn1_AV_readaddr(3),VMSTE_L4PHIAn1_AV_readaddr(2),VMSTE_L4PHIAn1_AV_readaddr(1),VMSTE_L4PHIAn1_AV_readaddr(0)),
        doutb     => VMSTE_L4PHIAn1_V_datatmp,
        enb_nent  => VMSTE_L4PHIAn1_enb_nent,
        addr_nent  => VMSTE_L4PHIAn1_V_addr_nent,
        dout_nent  => VMSTE_L4PHIAn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L4PHIAn1_enb_binmaska,
        addr_binmaska  => VMSTE_L4PHIAn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L4PHIAn1_V_binmaska,
        enb_binmaskb  => VMSTE_L4PHIAn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L4PHIAn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L4PHIAn1_V_binmaskb
      );

    VMSTE_L4PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L4PHIAn1_wea,
        addra     => VMSTE_L4PHIAn1_writeaddr,
        dina      => VMSTE_L4PHIAn1_din,
        wea_out       => VMSTE_L4PHIAn1_wea_delay,
        addra_out     => VMSTE_L4PHIAn1_writeaddr_delay,
        dina_out      => VMSTE_L4PHIAn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L4PHIAn1_start
      );

    VMSTE_L4PHIBn1_dataformat : entity work.vmstub17dout5
      port map (
        datain => VMSTE_L4PHIBn1_V_datatmp,
        dataout0 => VMSTE_L4PHIBn1_AV_dout(0),
        dataout1 => VMSTE_L4PHIBn1_AV_dout(1),
        dataout2 => VMSTE_L4PHIBn1_AV_dout(2),
        dataout3 => VMSTE_L4PHIBn1_AV_dout(3),
        dataout4 => VMSTE_L4PHIBn1_AV_dout(4)
      );

    VMSTE_L4PHIBn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L4PHIBn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L4PHIBn1_wea_delay,
        addra     => VMSTE_L4PHIBn1_writeaddr_delay,
        dina      => VMSTE_L4PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L4PHIBn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L4PHIBn1_AV_readaddr(4),VMSTE_L4PHIBn1_AV_readaddr(3),VMSTE_L4PHIBn1_AV_readaddr(2),VMSTE_L4PHIBn1_AV_readaddr(1),VMSTE_L4PHIBn1_AV_readaddr(0)),
        doutb     => VMSTE_L4PHIBn1_V_datatmp,
        enb_nent  => VMSTE_L4PHIBn1_enb_nent,
        addr_nent  => VMSTE_L4PHIBn1_V_addr_nent,
        dout_nent  => VMSTE_L4PHIBn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L4PHIBn1_enb_binmaska,
        addr_binmaska  => VMSTE_L4PHIBn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L4PHIBn1_V_binmaska,
        enb_binmaskb  => VMSTE_L4PHIBn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L4PHIBn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L4PHIBn1_V_binmaskb
      );

    VMSTE_L4PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L4PHIBn1_wea,
        addra     => VMSTE_L4PHIBn1_writeaddr,
        dina      => VMSTE_L4PHIBn1_din,
        wea_out       => VMSTE_L4PHIBn1_wea_delay,
        addra_out     => VMSTE_L4PHIBn1_writeaddr_delay,
        dina_out      => VMSTE_L4PHIBn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L4PHIBn1_start
      );

    VMSTE_L4PHICn1_dataformat : entity work.vmstub17dout5
      port map (
        datain => VMSTE_L4PHICn1_V_datatmp,
        dataout0 => VMSTE_L4PHICn1_AV_dout(0),
        dataout1 => VMSTE_L4PHICn1_AV_dout(1),
        dataout2 => VMSTE_L4PHICn1_AV_dout(2),
        dataout3 => VMSTE_L4PHICn1_AV_dout(3),
        dataout4 => VMSTE_L4PHICn1_AV_dout(4)
      );

    VMSTE_L4PHICn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L4PHICn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L4PHICn1_wea_delay,
        addra     => VMSTE_L4PHICn1_writeaddr_delay,
        dina      => VMSTE_L4PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L4PHICn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L4PHICn1_AV_readaddr(4),VMSTE_L4PHICn1_AV_readaddr(3),VMSTE_L4PHICn1_AV_readaddr(2),VMSTE_L4PHICn1_AV_readaddr(1),VMSTE_L4PHICn1_AV_readaddr(0)),
        doutb     => VMSTE_L4PHICn1_V_datatmp,
        enb_nent  => VMSTE_L4PHICn1_enb_nent,
        addr_nent  => VMSTE_L4PHICn1_V_addr_nent,
        dout_nent  => VMSTE_L4PHICn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L4PHICn1_enb_binmaska,
        addr_binmaska  => VMSTE_L4PHICn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L4PHICn1_V_binmaska,
        enb_binmaskb  => VMSTE_L4PHICn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L4PHICn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L4PHICn1_V_binmaskb
      );

    VMSTE_L4PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L4PHICn1_wea,
        addra     => VMSTE_L4PHICn1_writeaddr,
        dina      => VMSTE_L4PHICn1_din,
        wea_out       => VMSTE_L4PHICn1_wea_delay,
        addra_out     => VMSTE_L4PHICn1_writeaddr_delay,
        dina_out      => VMSTE_L4PHICn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L4PHICn1_start
      );

    VMSTE_L4PHIDn1_dataformat : entity work.vmstub17dout5
      port map (
        datain => VMSTE_L4PHIDn1_V_datatmp,
        dataout0 => VMSTE_L4PHIDn1_AV_dout(0),
        dataout1 => VMSTE_L4PHIDn1_AV_dout(1),
        dataout2 => VMSTE_L4PHIDn1_AV_dout(2),
        dataout3 => VMSTE_L4PHIDn1_AV_dout(3),
        dataout4 => VMSTE_L4PHIDn1_AV_dout(4)
      );

    VMSTE_L4PHIDn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L4PHIDn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 5
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L4PHIDn1_wea_delay,
        addra     => VMSTE_L4PHIDn1_writeaddr_delay,
        dina      => VMSTE_L4PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L4PHIDn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L4PHIDn1_AV_readaddr(4),VMSTE_L4PHIDn1_AV_readaddr(3),VMSTE_L4PHIDn1_AV_readaddr(2),VMSTE_L4PHIDn1_AV_readaddr(1),VMSTE_L4PHIDn1_AV_readaddr(0)),
        doutb     => VMSTE_L4PHIDn1_V_datatmp,
        enb_nent  => VMSTE_L4PHIDn1_enb_nent,
        addr_nent  => VMSTE_L4PHIDn1_V_addr_nent,
        dout_nent  => VMSTE_L4PHIDn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L4PHIDn1_enb_binmaska,
        addr_binmaska  => VMSTE_L4PHIDn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L4PHIDn1_V_binmaska,
        enb_binmaskb  => VMSTE_L4PHIDn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L4PHIDn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L4PHIDn1_V_binmaskb
      );

    VMSTE_L4PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L4PHIDn1_wea,
        addra     => VMSTE_L4PHIDn1_writeaddr,
        dina      => VMSTE_L4PHIDn1_din,
        wea_out       => VMSTE_L4PHIDn1_wea_delay,
        addra_out     => VMSTE_L4PHIDn1_writeaddr_delay,
        dina_out      => VMSTE_L4PHIDn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L4PHIDn1_start
      );

    VMSTE_L6PHIAn1_dataformat : entity work.vmstub17dout3
      port map (
        datain => VMSTE_L6PHIAn1_V_datatmp,
        dataout0 => VMSTE_L6PHIAn1_AV_dout(0),
        dataout1 => VMSTE_L6PHIAn1_AV_dout(1),
        dataout2 => VMSTE_L6PHIAn1_AV_dout(2)
      );

    VMSTE_L6PHIAn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L6PHIAn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L6PHIAn1_wea_delay,
        addra     => VMSTE_L6PHIAn1_writeaddr_delay,
        dina      => VMSTE_L6PHIAn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L6PHIAn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L6PHIAn1_AV_readaddr(2),VMSTE_L6PHIAn1_AV_readaddr(1),VMSTE_L6PHIAn1_AV_readaddr(0)),
        doutb     => VMSTE_L6PHIAn1_V_datatmp,
        enb_nent  => VMSTE_L6PHIAn1_enb_nent,
        addr_nent  => VMSTE_L6PHIAn1_V_addr_nent,
        dout_nent  => VMSTE_L6PHIAn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L6PHIAn1_enb_binmaska,
        addr_binmaska  => VMSTE_L6PHIAn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L6PHIAn1_V_binmaska,
        enb_binmaskb  => VMSTE_L6PHIAn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L6PHIAn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L6PHIAn1_V_binmaskb
      );

    VMSTE_L6PHIAn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L6PHIAn1_wea,
        addra     => VMSTE_L6PHIAn1_writeaddr,
        dina      => VMSTE_L6PHIAn1_din,
        wea_out       => VMSTE_L6PHIAn1_wea_delay,
        addra_out     => VMSTE_L6PHIAn1_writeaddr_delay,
        dina_out      => VMSTE_L6PHIAn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L6PHIAn1_start
      );

    VMSTE_L6PHIBn1_dataformat : entity work.vmstub17dout3
      port map (
        datain => VMSTE_L6PHIBn1_V_datatmp,
        dataout0 => VMSTE_L6PHIBn1_AV_dout(0),
        dataout1 => VMSTE_L6PHIBn1_AV_dout(1),
        dataout2 => VMSTE_L6PHIBn1_AV_dout(2)
      );

    VMSTE_L6PHIBn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L6PHIBn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L6PHIBn1_wea_delay,
        addra     => VMSTE_L6PHIBn1_writeaddr_delay,
        dina      => VMSTE_L6PHIBn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L6PHIBn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L6PHIBn1_AV_readaddr(2),VMSTE_L6PHIBn1_AV_readaddr(1),VMSTE_L6PHIBn1_AV_readaddr(0)),
        doutb     => VMSTE_L6PHIBn1_V_datatmp,
        enb_nent  => VMSTE_L6PHIBn1_enb_nent,
        addr_nent  => VMSTE_L6PHIBn1_V_addr_nent,
        dout_nent  => VMSTE_L6PHIBn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L6PHIBn1_enb_binmaska,
        addr_binmaska  => VMSTE_L6PHIBn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L6PHIBn1_V_binmaska,
        enb_binmaskb  => VMSTE_L6PHIBn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L6PHIBn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L6PHIBn1_V_binmaskb
      );

    VMSTE_L6PHIBn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L6PHIBn1_wea,
        addra     => VMSTE_L6PHIBn1_writeaddr,
        dina      => VMSTE_L6PHIBn1_din,
        wea_out       => VMSTE_L6PHIBn1_wea_delay,
        addra_out     => VMSTE_L6PHIBn1_writeaddr_delay,
        dina_out      => VMSTE_L6PHIBn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L6PHIBn1_start
      );

    VMSTE_L6PHICn1_dataformat : entity work.vmstub17dout3
      port map (
        datain => VMSTE_L6PHICn1_V_datatmp,
        dataout0 => VMSTE_L6PHICn1_AV_dout(0),
        dataout1 => VMSTE_L6PHICn1_AV_dout(1),
        dataout2 => VMSTE_L6PHICn1_AV_dout(2)
      );

    VMSTE_L6PHICn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L6PHICn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L6PHICn1_wea_delay,
        addra     => VMSTE_L6PHICn1_writeaddr_delay,
        dina      => VMSTE_L6PHICn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L6PHICn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L6PHICn1_AV_readaddr(2),VMSTE_L6PHICn1_AV_readaddr(1),VMSTE_L6PHICn1_AV_readaddr(0)),
        doutb     => VMSTE_L6PHICn1_V_datatmp,
        enb_nent  => VMSTE_L6PHICn1_enb_nent,
        addr_nent  => VMSTE_L6PHICn1_V_addr_nent,
        dout_nent  => VMSTE_L6PHICn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L6PHICn1_enb_binmaska,
        addr_binmaska  => VMSTE_L6PHICn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L6PHICn1_V_binmaska,
        enb_binmaskb  => VMSTE_L6PHICn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L6PHICn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L6PHICn1_V_binmaskb
      );

    VMSTE_L6PHICn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L6PHICn1_wea,
        addra     => VMSTE_L6PHICn1_writeaddr,
        dina      => VMSTE_L6PHICn1_din,
        wea_out       => VMSTE_L6PHICn1_wea_delay,
        addra_out     => VMSTE_L6PHICn1_writeaddr_delay,
        dina_out      => VMSTE_L6PHICn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L6PHICn1_start
      );

    VMSTE_L6PHIDn1_dataformat : entity work.vmstub17dout3
      port map (
        datain => VMSTE_L6PHIDn1_V_datatmp,
        dataout0 => VMSTE_L6PHIDn1_AV_dout(0),
        dataout1 => VMSTE_L6PHIDn1_AV_dout(1),
        dataout2 => VMSTE_L6PHIDn1_AV_dout(2)
      );

    VMSTE_L6PHIDn1 : entity work.tf_mem_bin
      generic map (
        RAM_WIDTH       => 17,
        NUM_PAGES       => 2,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "VMSTE_L6PHIDn1",
        ADDR_WIDTH      => 4,
        NUM_PHI_BINS    => 8,
        NUM_RZ_BINS     => 8,
        NUM_COPY        => 3
      )
      port map (
        clka      => clk,
        wea       => VMSTE_L6PHIDn1_wea_delay,
        addra     => VMSTE_L6PHIDn1_writeaddr_delay,
        dina      => VMSTE_L6PHIDn1_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        sync_nent => VMSTE_L6PHIDn1_start,
        enb       => (others => '1'),
        addrb     => (VMSTE_L6PHIDn1_AV_readaddr(2),VMSTE_L6PHIDn1_AV_readaddr(1),VMSTE_L6PHIDn1_AV_readaddr(0)),
        doutb     => VMSTE_L6PHIDn1_V_datatmp,
        enb_nent  => VMSTE_L6PHIDn1_enb_nent,
        addr_nent  => VMSTE_L6PHIDn1_V_addr_nent,
        dout_nent  => VMSTE_L6PHIDn1_AV_dout_nent,
        enb_binmaska  => VMSTE_L6PHIDn1_enb_binmaska,
        addr_binmaska  => VMSTE_L6PHIDn1_V_addr_binmaska,
        binmaska_o  => VMSTE_L6PHIDn1_V_binmaska,
        enb_binmaskb  => VMSTE_L6PHIDn1_enb_binmaskb,
        addr_binmaskb  => VMSTE_L6PHIDn1_V_addr_binmaskb,
        binmaskb_o  => VMSTE_L6PHIDn1_V_binmaskb
      );

    VMSTE_L6PHIDn1_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 2,
        RAM_DEPTH       => 2*PAGE_LENGTH_CM,
        RAM_WIDTH       => 17
      )
      port map (
        clk      => clk,
        wea       => VMSTE_L6PHIDn1_wea,
        addra     => VMSTE_L6PHIDn1_writeaddr,
        dina      => VMSTE_L6PHIDn1_din,
        wea_out       => VMSTE_L6PHIDn1_wea_delay,
        addra_out     => VMSTE_L6PHIDn1_writeaddr_delay,
        dina_out      => VMSTE_L6PHIDn1_din_delay,
        done       => VMR_done,
        start      => VMSTE_L6PHIDn1_start
      );

    TPARL1L2ABC_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1L2ABC_bx,
        bx_vld => TPARL1L2ABC_bx_vld
      );

--    MERGE_STREAM_TPARL1L2ABC : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 3,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1L2ABC_bx,
--        bx_in_vld => TPARL1L2ABC_bx_vld,
--        rst => '0',
--        clk => clk,
--        bx_out => TP_bx_out_merged,
--        merged_dout => MPAR_L1L2ABC_stream_V_dout,
--        din0=>TPAR_L1L2A_V_dout,
--        din1=>TPAR_L1L2B_V_dout,
--        din2=>TPAR_L1L2C_V_dout,
--        din3=>TPAR_L1L2A_V_dout,
--        nent0=>TPAR_L1L2A_AV_dout_nent,
--        nent1=>TPAR_L1L2B_AV_dout_nent,
--        nent2=>TPAR_L1L2C_AV_dout_nent,
--        nent3=>TPAR_L1L2A_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1L2A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L1L2B_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_L1L2C_V_readaddr
--      );

    TPAR_L1L2A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2A_wea_delay,
        addra     => TPAR_L1L2A_writeaddr_delay,
        dina      => TPAR_L1L2A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2A_V_readaddr,
        doutb     => TPAR_L1L2A_V_dout,
        sync_nent => TPAR_L1L2A_start,
        nent_o    => TPAR_L1L2A_AV_dout_nent
      );

    TPAR_L1L2A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2A_wea,
        addra     => TPAR_L1L2A_writeaddr,
        dina      => TPAR_L1L2A_din,
        wea_out       => TPAR_L1L2A_wea_delay,
        addra_out     => TPAR_L1L2A_writeaddr_delay,
        dina_out      => TPAR_L1L2A_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2A_start
      );

    TPAR_L1L2B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2B_wea_delay,
        addra     => TPAR_L1L2B_writeaddr_delay,
        dina      => TPAR_L1L2B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2B_V_readaddr,
        doutb     => TPAR_L1L2B_V_dout,
        sync_nent => TPAR_L1L2B_start,
        nent_o    => TPAR_L1L2B_AV_dout_nent
      );

    TPAR_L1L2B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2B_wea,
        addra     => TPAR_L1L2B_writeaddr,
        dina      => TPAR_L1L2B_din,
        wea_out       => TPAR_L1L2B_wea_delay,
        addra_out     => TPAR_L1L2B_writeaddr_delay,
        dina_out      => TPAR_L1L2B_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2B_start
      );

    TPAR_L1L2C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2C_wea_delay,
        addra     => TPAR_L1L2C_writeaddr_delay,
        dina      => TPAR_L1L2C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2C_V_readaddr,
        doutb     => TPAR_L1L2C_V_dout,
        sync_nent => TPAR_L1L2C_start,
        nent_o    => TPAR_L1L2C_AV_dout_nent
      );

    TPAR_L1L2C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2C_wea,
        addra     => TPAR_L1L2C_writeaddr,
        dina      => TPAR_L1L2C_din,
        wea_out       => TPAR_L1L2C_wea_delay,
        addra_out     => TPAR_L1L2C_writeaddr_delay,
        dina_out      => TPAR_L1L2C_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2C_start
      );

    TPARL1L2DE_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1L2DE_bx,
        bx_vld => TPARL1L2DE_bx_vld
      );

--    MERGE_STREAM_TPARL1L2DE : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 2,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1L2DE_bx,
--        bx_in_vld => TPARL1L2DE_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L1L2DE_stream_V_dout,
--        din0=>TPAR_L1L2D_V_dout,
--        din1=>TPAR_L1L2E_V_dout,
--        din2=>TPAR_L1L2D_V_dout,
--        din3=>TPAR_L1L2E_V_dout,
--        nent0=>TPAR_L1L2D_AV_dout_nent,
--        nent1=>TPAR_L1L2E_AV_dout_nent,
--        nent2=>TPAR_L1L2D_AV_dout_nent,
--        nent3=>TPAR_L1L2E_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1L2D_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L1L2E_V_readaddr
--      );

    TPAR_L1L2D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2D_wea_delay,
        addra     => TPAR_L1L2D_writeaddr_delay,
        dina      => TPAR_L1L2D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2D_V_readaddr,
        doutb     => TPAR_L1L2D_V_dout,
        sync_nent => TPAR_L1L2D_start,
        nent_o    => TPAR_L1L2D_AV_dout_nent
      );

    TPAR_L1L2D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2D_wea,
        addra     => TPAR_L1L2D_writeaddr,
        dina      => TPAR_L1L2D_din,
        wea_out       => TPAR_L1L2D_wea_delay,
        addra_out     => TPAR_L1L2D_writeaddr_delay,
        dina_out      => TPAR_L1L2D_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2D_start
      );

    TPAR_L1L2E : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2E",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2E_wea_delay,
        addra     => TPAR_L1L2E_writeaddr_delay,
        dina      => TPAR_L1L2E_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2E_V_readaddr,
        doutb     => TPAR_L1L2E_V_dout,
        sync_nent => TPAR_L1L2E_start,
        nent_o    => TPAR_L1L2E_AV_dout_nent
      );

    TPAR_L1L2E_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2E_wea,
        addra     => TPAR_L1L2E_writeaddr,
        dina      => TPAR_L1L2E_din,
        wea_out       => TPAR_L1L2E_wea_delay,
        addra_out     => TPAR_L1L2E_writeaddr_delay,
        dina_out      => TPAR_L1L2E_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2E_start
      );

    TPARL1L2F_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1L2F_bx,
        bx_vld => TPARL1L2F_bx_vld
      );

--    MERGE_STREAM_TPARL1L2F : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1L2F_bx,
--        bx_in_vld => TPARL1L2F_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L1L2F_stream_V_dout,
--        din0=>TPAR_L1L2F_V_dout,
--        din1=>TPAR_L1L2F_V_dout,
--        din2=>TPAR_L1L2F_V_dout,
--        din3=>TPAR_L1L2F_V_dout,
--        nent0=>TPAR_L1L2F_AV_dout_nent,
--        nent1=>TPAR_L1L2F_AV_dout_nent,
--        nent2=>TPAR_L1L2F_AV_dout_nent,
--        nent3=>TPAR_L1L2F_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1L2F_V_readaddr
--      );

    TPAR_L1L2F : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2F",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2F_wea_delay,
        addra     => TPAR_L1L2F_writeaddr_delay,
        dina      => TPAR_L1L2F_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2F_V_readaddr,
        doutb     => TPAR_L1L2F_V_dout,
        sync_nent => TPAR_L1L2F_start,
        nent_o    => TPAR_L1L2F_AV_dout_nent
      );

    TPAR_L1L2F_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2F_wea,
        addra     => TPAR_L1L2F_writeaddr,
        dina      => TPAR_L1L2F_din,
        wea_out       => TPAR_L1L2F_wea_delay,
        addra_out     => TPAR_L1L2F_writeaddr_delay,
        dina_out      => TPAR_L1L2F_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2F_start
      );

    TPARL1L2G_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1L2G_bx,
        bx_vld => TPARL1L2G_bx_vld
      );

--    MERGE_STREAM_TPARL1L2G : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 1,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1L2G_bx,
--        bx_in_vld => TPARL1L2G_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L1L2G_stream_V_dout,
--        din0=>TPAR_L1L2G_V_dout,
--        din1=>TPAR_L1L2G_V_dout,
--        din2=>TPAR_L1L2G_V_dout,
--        din3=>TPAR_L1L2G_V_dout,
--        nent0=>TPAR_L1L2G_AV_dout_nent,
--        nent1=>TPAR_L1L2G_AV_dout_nent,
--        nent2=>TPAR_L1L2G_AV_dout_nent,
--        nent3=>TPAR_L1L2G_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1L2G_V_readaddr
--      );

    TPAR_L1L2G : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2G",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2G_wea_delay,
        addra     => TPAR_L1L2G_writeaddr_delay,
        dina      => TPAR_L1L2G_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2G_V_readaddr,
        doutb     => TPAR_L1L2G_V_dout,
        sync_nent => TPAR_L1L2G_start,
        nent_o    => TPAR_L1L2G_AV_dout_nent
      );

    TPAR_L1L2G_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2G_wea,
        addra     => TPAR_L1L2G_writeaddr,
        dina      => TPAR_L1L2G_din,
        wea_out       => TPAR_L1L2G_wea_delay,
        addra_out     => TPAR_L1L2G_writeaddr_delay,
        dina_out      => TPAR_L1L2G_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2G_start
      );

    TPARL1L2HI_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1L2HI_bx,
        bx_vld => TPARL1L2HI_bx_vld
      );

--    MERGE_STREAM_TPARL1L2HI : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 2,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1L2HI_bx,
--        bx_in_vld => TPARL1L2HI_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L1L2HI_stream_V_dout,
--        din0=>TPAR_L1L2H_V_dout,
--        din1=>TPAR_L1L2I_V_dout,
--        din2=>TPAR_L1L2H_V_dout,
--        din3=>TPAR_L1L2I_V_dout,
--        nent0=>TPAR_L1L2H_AV_dout_nent,
--        nent1=>TPAR_L1L2I_AV_dout_nent,
--        nent2=>TPAR_L1L2H_AV_dout_nent,
--        nent3=>TPAR_L1L2I_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1L2H_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L1L2I_V_readaddr
--      );

    TPAR_L1L2H : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2H",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2H_wea_delay,
        addra     => TPAR_L1L2H_writeaddr_delay,
        dina      => TPAR_L1L2H_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2H_V_readaddr,
        doutb     => TPAR_L1L2H_V_dout,
        sync_nent => TPAR_L1L2H_start,
        nent_o    => TPAR_L1L2H_AV_dout_nent
      );

    TPAR_L1L2H_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2H_wea,
        addra     => TPAR_L1L2H_writeaddr,
        dina      => TPAR_L1L2H_din,
        wea_out       => TPAR_L1L2H_wea_delay,
        addra_out     => TPAR_L1L2H_writeaddr_delay,
        dina_out      => TPAR_L1L2H_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2H_start
      );

    TPAR_L1L2I : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2I",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2I_wea_delay,
        addra     => TPAR_L1L2I_writeaddr_delay,
        dina      => TPAR_L1L2I_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2I_V_readaddr,
        doutb     => TPAR_L1L2I_V_dout,
        sync_nent => TPAR_L1L2I_start,
        nent_o    => TPAR_L1L2I_AV_dout_nent
      );

    TPAR_L1L2I_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2I_wea,
        addra     => TPAR_L1L2I_writeaddr,
        dina      => TPAR_L1L2I_din,
        wea_out       => TPAR_L1L2I_wea_delay,
        addra_out     => TPAR_L1L2I_writeaddr_delay,
        dina_out      => TPAR_L1L2I_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2I_start
      );

    TPARL1L2JKL_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1L2JKL_bx,
        bx_vld => TPARL1L2JKL_bx_vld
      );

--    MERGE_STREAM_TPARL1L2JKL : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 3,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1L2JKL_bx,
--        bx_in_vld => TPARL1L2JKL_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L1L2JKL_stream_V_dout,
--        din0=>TPAR_L1L2J_V_dout,
--        din1=>TPAR_L1L2K_V_dout,
--        din2=>TPAR_L1L2L_V_dout,
--        din3=>TPAR_L1L2J_V_dout,
--        nent0=>TPAR_L1L2J_AV_dout_nent,
--        nent1=>TPAR_L1L2K_AV_dout_nent,
--        nent2=>TPAR_L1L2L_AV_dout_nent,
--        nent3=>TPAR_L1L2J_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1L2J_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L1L2K_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_L1L2L_V_readaddr
--      );

    TPAR_L1L2J : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2J",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2J_wea_delay,
        addra     => TPAR_L1L2J_writeaddr_delay,
        dina      => TPAR_L1L2J_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2J_V_readaddr,
        doutb     => TPAR_L1L2J_V_dout,
        sync_nent => TPAR_L1L2J_start,
        nent_o    => TPAR_L1L2J_AV_dout_nent
      );

    TPAR_L1L2J_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2J_wea,
        addra     => TPAR_L1L2J_writeaddr,
        dina      => TPAR_L1L2J_din,
        wea_out       => TPAR_L1L2J_wea_delay,
        addra_out     => TPAR_L1L2J_writeaddr_delay,
        dina_out      => TPAR_L1L2J_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2J_start
      );

    TPAR_L1L2K : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2K",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2K_wea_delay,
        addra     => TPAR_L1L2K_writeaddr_delay,
        dina      => TPAR_L1L2K_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2K_V_readaddr,
        doutb     => TPAR_L1L2K_V_dout,
        sync_nent => TPAR_L1L2K_start,
        nent_o    => TPAR_L1L2K_AV_dout_nent
      );

    TPAR_L1L2K_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2K_wea,
        addra     => TPAR_L1L2K_writeaddr,
        dina      => TPAR_L1L2K_din,
        wea_out       => TPAR_L1L2K_wea_delay,
        addra_out     => TPAR_L1L2K_writeaddr_delay,
        dina_out      => TPAR_L1L2K_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2K_start
      );

    TPAR_L1L2L : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1L2L",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1L2L_wea_delay,
        addra     => TPAR_L1L2L_writeaddr_delay,
        dina      => TPAR_L1L2L_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1L2L_V_readaddr,
        doutb     => TPAR_L1L2L_V_dout,
        sync_nent => TPAR_L1L2L_start,
        nent_o    => TPAR_L1L2L_AV_dout_nent
      );

    TPAR_L1L2L_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1L2L_wea,
        addra     => TPAR_L1L2L_writeaddr,
        dina      => TPAR_L1L2L_din,
        wea_out       => TPAR_L1L2L_wea_delay,
        addra_out     => TPAR_L1L2L_writeaddr_delay,
        dina_out      => TPAR_L1L2L_din_delay,
        done       => TP_done,
        start      => TPAR_L1L2L_start
      );

    TPARL2L3ABCD_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL2L3ABCD_bx,
        bx_vld => TPARL2L3ABCD_bx_vld
      );

--    MERGE_STREAM_TPARL2L3ABCD : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 4,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL2L3ABCD_bx,
--        bx_in_vld => TPARL2L3ABCD_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L2L3ABCD_stream_V_dout,
--        din0=>TPAR_L2L3A_V_dout,
--        din1=>TPAR_L2L3B_V_dout,
--        din2=>TPAR_L2L3C_V_dout,
--        din3=>TPAR_L2L3D_V_dout,
--        nent0=>TPAR_L2L3A_AV_dout_nent,
--        nent1=>TPAR_L2L3B_AV_dout_nent,
--        nent2=>TPAR_L2L3C_AV_dout_nent,
--        nent3=>TPAR_L2L3D_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L2L3A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L2L3B_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_L2L3C_V_readaddr,
--        addr_arr(39 downto 30)=>TPAR_L2L3D_V_readaddr
--      );

    TPAR_L2L3A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2L3A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2L3A_wea_delay,
        addra     => TPAR_L2L3A_writeaddr_delay,
        dina      => TPAR_L2L3A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2L3A_V_readaddr,
        doutb     => TPAR_L2L3A_V_dout,
        sync_nent => TPAR_L2L3A_start,
        nent_o    => TPAR_L2L3A_AV_dout_nent
      );

    TPAR_L2L3A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2L3A_wea,
        addra     => TPAR_L2L3A_writeaddr,
        dina      => TPAR_L2L3A_din,
        wea_out       => TPAR_L2L3A_wea_delay,
        addra_out     => TPAR_L2L3A_writeaddr_delay,
        dina_out      => TPAR_L2L3A_din_delay,
        done       => TP_done,
        start      => TPAR_L2L3A_start
      );

    TPAR_L2L3B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2L3B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2L3B_wea_delay,
        addra     => TPAR_L2L3B_writeaddr_delay,
        dina      => TPAR_L2L3B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2L3B_V_readaddr,
        doutb     => TPAR_L2L3B_V_dout,
        sync_nent => TPAR_L2L3B_start,
        nent_o    => TPAR_L2L3B_AV_dout_nent
      );

    TPAR_L2L3B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2L3B_wea,
        addra     => TPAR_L2L3B_writeaddr,
        dina      => TPAR_L2L3B_din,
        wea_out       => TPAR_L2L3B_wea_delay,
        addra_out     => TPAR_L2L3B_writeaddr_delay,
        dina_out      => TPAR_L2L3B_din_delay,
        done       => TP_done,
        start      => TPAR_L2L3B_start
      );

    TPAR_L2L3C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2L3C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2L3C_wea_delay,
        addra     => TPAR_L2L3C_writeaddr_delay,
        dina      => TPAR_L2L3C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2L3C_V_readaddr,
        doutb     => TPAR_L2L3C_V_dout,
        sync_nent => TPAR_L2L3C_start,
        nent_o    => TPAR_L2L3C_AV_dout_nent
      );

    TPAR_L2L3C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2L3C_wea,
        addra     => TPAR_L2L3C_writeaddr,
        dina      => TPAR_L2L3C_din,
        wea_out       => TPAR_L2L3C_wea_delay,
        addra_out     => TPAR_L2L3C_writeaddr_delay,
        dina_out      => TPAR_L2L3C_din_delay,
        done       => TP_done,
        start      => TPAR_L2L3C_start
      );

    TPAR_L2L3D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2L3D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2L3D_wea_delay,
        addra     => TPAR_L2L3D_writeaddr_delay,
        dina      => TPAR_L2L3D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2L3D_V_readaddr,
        doutb     => TPAR_L2L3D_V_dout,
        sync_nent => TPAR_L2L3D_start,
        nent_o    => TPAR_L2L3D_AV_dout_nent
      );

    TPAR_L2L3D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2L3D_wea,
        addra     => TPAR_L2L3D_writeaddr,
        dina      => TPAR_L2L3D_din,
        wea_out       => TPAR_L2L3D_wea_delay,
        addra_out     => TPAR_L2L3D_writeaddr_delay,
        dina_out      => TPAR_L2L3D_din_delay,
        done       => TP_done,
        start      => TPAR_L2L3D_start
      );

    TPARL3L4AB_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL3L4AB_bx,
        bx_vld => TPARL3L4AB_bx_vld
      );

--    MERGE_STREAM_TPARL3L4AB : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 2,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL3L4AB_bx,
--        bx_in_vld => TPARL3L4AB_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L3L4AB_stream_V_dout,
--        din0=>TPAR_L3L4A_V_dout,
--        din1=>TPAR_L3L4B_V_dout,
--        din2=>TPAR_L3L4A_V_dout,
--        din3=>TPAR_L3L4B_V_dout,
--        nent0=>TPAR_L3L4A_AV_dout_nent,
--        nent1=>TPAR_L3L4B_AV_dout_nent,
--        nent2=>TPAR_L3L4A_AV_dout_nent,
--        nent3=>TPAR_L3L4B_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L3L4A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L3L4B_V_readaddr
--      );

    TPAR_L3L4A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L3L4A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L3L4A_wea_delay,
        addra     => TPAR_L3L4A_writeaddr_delay,
        dina      => TPAR_L3L4A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L3L4A_V_readaddr,
        doutb     => TPAR_L3L4A_V_dout,
        sync_nent => TPAR_L3L4A_start,
        nent_o    => TPAR_L3L4A_AV_dout_nent
      );

    TPAR_L3L4A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L3L4A_wea,
        addra     => TPAR_L3L4A_writeaddr,
        dina      => TPAR_L3L4A_din,
        wea_out       => TPAR_L3L4A_wea_delay,
        addra_out     => TPAR_L3L4A_writeaddr_delay,
        dina_out      => TPAR_L3L4A_din_delay,
        done       => TP_done,
        start      => TPAR_L3L4A_start
      );

    TPAR_L3L4B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L3L4B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L3L4B_wea_delay,
        addra     => TPAR_L3L4B_writeaddr_delay,
        dina      => TPAR_L3L4B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L3L4B_V_readaddr,
        doutb     => TPAR_L3L4B_V_dout,
        sync_nent => TPAR_L3L4B_start,
        nent_o    => TPAR_L3L4B_AV_dout_nent
      );

    TPAR_L3L4B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L3L4B_wea,
        addra     => TPAR_L3L4B_writeaddr,
        dina      => TPAR_L3L4B_din,
        wea_out       => TPAR_L3L4B_wea_delay,
        addra_out     => TPAR_L3L4B_writeaddr_delay,
        dina_out      => TPAR_L3L4B_din_delay,
        done       => TP_done,
        start      => TPAR_L3L4B_start
      );

    TPARL3L4CD_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL3L4CD_bx,
        bx_vld => TPARL3L4CD_bx_vld
      );

--    MERGE_STREAM_TPARL3L4CD : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 2,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL3L4CD_bx,
--        bx_in_vld => TPARL3L4CD_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L3L4CD_stream_V_dout,
--        din0=>TPAR_L3L4C_V_dout,
--        din1=>TPAR_L3L4D_V_dout,
--        din2=>TPAR_L3L4C_V_dout,
--        din3=>TPAR_L3L4D_V_dout,
--        nent0=>TPAR_L3L4C_AV_dout_nent,
--        nent1=>TPAR_L3L4D_AV_dout_nent,
--        nent2=>TPAR_L3L4C_AV_dout_nent,
--        nent3=>TPAR_L3L4D_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L3L4C_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L3L4D_V_readaddr
--      );

    TPAR_L3L4C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L3L4C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L3L4C_wea_delay,
        addra     => TPAR_L3L4C_writeaddr_delay,
        dina      => TPAR_L3L4C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L3L4C_V_readaddr,
        doutb     => TPAR_L3L4C_V_dout,
        sync_nent => TPAR_L3L4C_start,
        nent_o    => TPAR_L3L4C_AV_dout_nent
      );

    TPAR_L3L4C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L3L4C_wea,
        addra     => TPAR_L3L4C_writeaddr,
        dina      => TPAR_L3L4C_din,
        wea_out       => TPAR_L3L4C_wea_delay,
        addra_out     => TPAR_L3L4C_writeaddr_delay,
        dina_out      => TPAR_L3L4C_din_delay,
        done       => TP_done,
        start      => TPAR_L3L4C_start
      );

    TPAR_L3L4D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L3L4D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L3L4D_wea_delay,
        addra     => TPAR_L3L4D_writeaddr_delay,
        dina      => TPAR_L3L4D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L3L4D_V_readaddr,
        doutb     => TPAR_L3L4D_V_dout,
        sync_nent => TPAR_L3L4D_start,
        nent_o    => TPAR_L3L4D_AV_dout_nent
      );

    TPAR_L3L4D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L3L4D_wea,
        addra     => TPAR_L3L4D_writeaddr,
        dina      => TPAR_L3L4D_din,
        wea_out       => TPAR_L3L4D_wea_delay,
        addra_out     => TPAR_L3L4D_writeaddr_delay,
        dina_out      => TPAR_L3L4D_din_delay,
        done       => TP_done,
        start      => TPAR_L3L4D_start
      );

    TPARL5L6ABCD_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL5L6ABCD_bx,
        bx_vld => TPARL5L6ABCD_bx_vld
      );

--    MERGE_STREAM_TPARL5L6ABCD : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 4,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL5L6ABCD_bx,
--        bx_in_vld => TPARL5L6ABCD_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L5L6ABCD_stream_V_dout,
--        din0=>TPAR_L5L6A_V_dout,
--        din1=>TPAR_L5L6B_V_dout,
--        din2=>TPAR_L5L6C_V_dout,
--        din3=>TPAR_L5L6D_V_dout,
--        nent0=>TPAR_L5L6A_AV_dout_nent,
--        nent1=>TPAR_L5L6B_AV_dout_nent,
--        nent2=>TPAR_L5L6C_AV_dout_nent,
--        nent3=>TPAR_L5L6D_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L5L6A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L5L6B_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_L5L6C_V_readaddr,
--        addr_arr(39 downto 30)=>TPAR_L5L6D_V_readaddr
--      );

    TPAR_L5L6A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L5L6A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L5L6A_wea_delay,
        addra     => TPAR_L5L6A_writeaddr_delay,
        dina      => TPAR_L5L6A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L5L6A_V_readaddr,
        doutb     => TPAR_L5L6A_V_dout,
        sync_nent => TPAR_L5L6A_start,
        nent_o    => TPAR_L5L6A_AV_dout_nent
      );

    TPAR_L5L6A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L5L6A_wea,
        addra     => TPAR_L5L6A_writeaddr,
        dina      => TPAR_L5L6A_din,
        wea_out       => TPAR_L5L6A_wea_delay,
        addra_out     => TPAR_L5L6A_writeaddr_delay,
        dina_out      => TPAR_L5L6A_din_delay,
        done       => TP_done,
        start      => TPAR_L5L6A_start
      );

    TPAR_L5L6B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L5L6B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L5L6B_wea_delay,
        addra     => TPAR_L5L6B_writeaddr_delay,
        dina      => TPAR_L5L6B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L5L6B_V_readaddr,
        doutb     => TPAR_L5L6B_V_dout,
        sync_nent => TPAR_L5L6B_start,
        nent_o    => TPAR_L5L6B_AV_dout_nent
      );

    TPAR_L5L6B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L5L6B_wea,
        addra     => TPAR_L5L6B_writeaddr,
        dina      => TPAR_L5L6B_din,
        wea_out       => TPAR_L5L6B_wea_delay,
        addra_out     => TPAR_L5L6B_writeaddr_delay,
        dina_out      => TPAR_L5L6B_din_delay,
        done       => TP_done,
        start      => TPAR_L5L6B_start
      );

    TPAR_L5L6C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L5L6C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L5L6C_wea_delay,
        addra     => TPAR_L5L6C_writeaddr_delay,
        dina      => TPAR_L5L6C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L5L6C_V_readaddr,
        doutb     => TPAR_L5L6C_V_dout,
        sync_nent => TPAR_L5L6C_start,
        nent_o    => TPAR_L5L6C_AV_dout_nent
      );

    TPAR_L5L6C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L5L6C_wea,
        addra     => TPAR_L5L6C_writeaddr,
        dina      => TPAR_L5L6C_din,
        wea_out       => TPAR_L5L6C_wea_delay,
        addra_out     => TPAR_L5L6C_writeaddr_delay,
        dina_out      => TPAR_L5L6C_din_delay,
        done       => TP_done,
        start      => TPAR_L5L6C_start
      );

    TPAR_L5L6D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L5L6D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L5L6D_wea_delay,
        addra     => TPAR_L5L6D_writeaddr_delay,
        dina      => TPAR_L5L6D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L5L6D_V_readaddr,
        doutb     => TPAR_L5L6D_V_dout,
        sync_nent => TPAR_L5L6D_start,
        nent_o    => TPAR_L5L6D_AV_dout_nent
      );

    TPAR_L5L6D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L5L6D_wea,
        addra     => TPAR_L5L6D_writeaddr,
        dina      => TPAR_L5L6D_din,
        wea_out       => TPAR_L5L6D_wea_delay,
        addra_out     => TPAR_L5L6D_writeaddr_delay,
        dina_out      => TPAR_L5L6D_din_delay,
        done       => TP_done,
        start      => TPAR_L5L6D_start
      );

    TPARD1D2ABCD_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARD1D2ABCD_bx,
        bx_vld => TPARD1D2ABCD_bx_vld
      );

--    MERGE_STREAM_TPARD1D2ABCD : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 4,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARD1D2ABCD_bx,
--        bx_in_vld => TPARD1D2ABCD_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_D1D2ABCD_stream_V_dout,
--        din0=>TPAR_D1D2A_V_dout,
--        din1=>TPAR_D1D2B_V_dout,
--        din2=>TPAR_D1D2C_V_dout,
--        din3=>TPAR_D1D2D_V_dout,
--        nent0=>TPAR_D1D2A_AV_dout_nent,
--        nent1=>TPAR_D1D2B_AV_dout_nent,
--        nent2=>TPAR_D1D2C_AV_dout_nent,
--        nent3=>TPAR_D1D2D_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_D1D2A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_D1D2B_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_D1D2C_V_readaddr,
--        addr_arr(39 downto 30)=>TPAR_D1D2D_V_readaddr
--      );

    TPAR_D1D2A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D1D2A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D1D2A_wea_delay,
        addra     => TPAR_D1D2A_writeaddr_delay,
        dina      => TPAR_D1D2A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D1D2A_V_readaddr,
        doutb     => TPAR_D1D2A_V_dout,
        sync_nent => TPAR_D1D2A_start,
        nent_o    => TPAR_D1D2A_AV_dout_nent
      );

    TPAR_D1D2A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D1D2A_wea,
        addra     => TPAR_D1D2A_writeaddr,
        dina      => TPAR_D1D2A_din,
        wea_out       => TPAR_D1D2A_wea_delay,
        addra_out     => TPAR_D1D2A_writeaddr_delay,
        dina_out      => TPAR_D1D2A_din_delay,
        done       => TP_done,
        start      => TPAR_D1D2A_start
      );

    TPAR_D1D2B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D1D2B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D1D2B_wea_delay,
        addra     => TPAR_D1D2B_writeaddr_delay,
        dina      => TPAR_D1D2B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D1D2B_V_readaddr,
        doutb     => TPAR_D1D2B_V_dout,
        sync_nent => TPAR_D1D2B_start,
        nent_o    => TPAR_D1D2B_AV_dout_nent
      );

    TPAR_D1D2B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D1D2B_wea,
        addra     => TPAR_D1D2B_writeaddr,
        dina      => TPAR_D1D2B_din,
        wea_out       => TPAR_D1D2B_wea_delay,
        addra_out     => TPAR_D1D2B_writeaddr_delay,
        dina_out      => TPAR_D1D2B_din_delay,
        done       => TP_done,
        start      => TPAR_D1D2B_start
      );

    TPAR_D1D2C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D1D2C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D1D2C_wea_delay,
        addra     => TPAR_D1D2C_writeaddr_delay,
        dina      => TPAR_D1D2C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D1D2C_V_readaddr,
        doutb     => TPAR_D1D2C_V_dout,
        sync_nent => TPAR_D1D2C_start,
        nent_o    => TPAR_D1D2C_AV_dout_nent
      );

    TPAR_D1D2C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D1D2C_wea,
        addra     => TPAR_D1D2C_writeaddr,
        dina      => TPAR_D1D2C_din,
        wea_out       => TPAR_D1D2C_wea_delay,
        addra_out     => TPAR_D1D2C_writeaddr_delay,
        dina_out      => TPAR_D1D2C_din_delay,
        done       => TP_done,
        start      => TPAR_D1D2C_start
      );

    TPAR_D1D2D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D1D2D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D1D2D_wea_delay,
        addra     => TPAR_D1D2D_writeaddr_delay,
        dina      => TPAR_D1D2D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D1D2D_V_readaddr,
        doutb     => TPAR_D1D2D_V_dout,
        sync_nent => TPAR_D1D2D_start,
        nent_o    => TPAR_D1D2D_AV_dout_nent
      );

    TPAR_D1D2D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D1D2D_wea,
        addra     => TPAR_D1D2D_writeaddr,
        dina      => TPAR_D1D2D_din,
        wea_out       => TPAR_D1D2D_wea_delay,
        addra_out     => TPAR_D1D2D_writeaddr_delay,
        dina_out      => TPAR_D1D2D_din_delay,
        done       => TP_done,
        start      => TPAR_D1D2D_start
      );

    TPARD3D4ABCD_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARD3D4ABCD_bx,
        bx_vld => TPARD3D4ABCD_bx_vld
      );

--    MERGE_STREAM_TPARD3D4ABCD : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 4,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARD3D4ABCD_bx,
--        bx_in_vld => TPARD3D4ABCD_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_D3D4ABCD_stream_V_dout,
--        din0=>TPAR_D3D4A_V_dout,
--        din1=>TPAR_D3D4B_V_dout,
--        din2=>TPAR_D3D4C_V_dout,
--        din3=>TPAR_D3D4D_V_dout,
--        nent0=>TPAR_D3D4A_AV_dout_nent,
--        nent1=>TPAR_D3D4B_AV_dout_nent,
--        nent2=>TPAR_D3D4C_AV_dout_nent,
--        nent3=>TPAR_D3D4D_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_D3D4A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_D3D4B_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_D3D4C_V_readaddr,
--        addr_arr(39 downto 30)=>TPAR_D3D4D_V_readaddr
--      );

    TPAR_D3D4A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D3D4A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D3D4A_wea_delay,
        addra     => TPAR_D3D4A_writeaddr_delay,
        dina      => TPAR_D3D4A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D3D4A_V_readaddr,
        doutb     => TPAR_D3D4A_V_dout,
        sync_nent => TPAR_D3D4A_start,
        nent_o    => TPAR_D3D4A_AV_dout_nent
      );

    TPAR_D3D4A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D3D4A_wea,
        addra     => TPAR_D3D4A_writeaddr,
        dina      => TPAR_D3D4A_din,
        wea_out       => TPAR_D3D4A_wea_delay,
        addra_out     => TPAR_D3D4A_writeaddr_delay,
        dina_out      => TPAR_D3D4A_din_delay,
        done       => TP_done,
        start      => TPAR_D3D4A_start
      );

    TPAR_D3D4B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D3D4B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D3D4B_wea_delay,
        addra     => TPAR_D3D4B_writeaddr_delay,
        dina      => TPAR_D3D4B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D3D4B_V_readaddr,
        doutb     => TPAR_D3D4B_V_dout,
        sync_nent => TPAR_D3D4B_start,
        nent_o    => TPAR_D3D4B_AV_dout_nent
      );

    TPAR_D3D4B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D3D4B_wea,
        addra     => TPAR_D3D4B_writeaddr,
        dina      => TPAR_D3D4B_din,
        wea_out       => TPAR_D3D4B_wea_delay,
        addra_out     => TPAR_D3D4B_writeaddr_delay,
        dina_out      => TPAR_D3D4B_din_delay,
        done       => TP_done,
        start      => TPAR_D3D4B_start
      );

    TPAR_D3D4C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D3D4C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D3D4C_wea_delay,
        addra     => TPAR_D3D4C_writeaddr_delay,
        dina      => TPAR_D3D4C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D3D4C_V_readaddr,
        doutb     => TPAR_D3D4C_V_dout,
        sync_nent => TPAR_D3D4C_start,
        nent_o    => TPAR_D3D4C_AV_dout_nent
      );

    TPAR_D3D4C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D3D4C_wea,
        addra     => TPAR_D3D4C_writeaddr,
        dina      => TPAR_D3D4C_din,
        wea_out       => TPAR_D3D4C_wea_delay,
        addra_out     => TPAR_D3D4C_writeaddr_delay,
        dina_out      => TPAR_D3D4C_din_delay,
        done       => TP_done,
        start      => TPAR_D3D4C_start
      );

    TPAR_D3D4D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_D3D4D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_D3D4D_wea_delay,
        addra     => TPAR_D3D4D_writeaddr_delay,
        dina      => TPAR_D3D4D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_D3D4D_V_readaddr,
        doutb     => TPAR_D3D4D_V_dout,
        sync_nent => TPAR_D3D4D_start,
        nent_o    => TPAR_D3D4D_AV_dout_nent
      );

    TPAR_D3D4D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_D3D4D_wea,
        addra     => TPAR_D3D4D_writeaddr,
        dina      => TPAR_D3D4D_din,
        wea_out       => TPAR_D3D4D_wea_delay,
        addra_out     => TPAR_D3D4D_writeaddr_delay,
        dina_out      => TPAR_D3D4D_din_delay,
        done       => TP_done,
        start      => TPAR_D3D4D_start
      );

    TPARL1D1ABCD_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1D1ABCD_bx,
        bx_vld => TPARL1D1ABCD_bx_vld
      );

--    MERGE_STREAM_TPARL1D1ABCD : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 4,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1D1ABCD_bx,
--        bx_in_vld => TPARL1D1ABCD_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L1D1ABCD_stream_V_dout,
--        din0=>TPAR_L1D1A_V_dout,
--        din1=>TPAR_L1D1B_V_dout,
--        din2=>TPAR_L1D1C_V_dout,
--        din3=>TPAR_L1D1D_V_dout,
--        nent0=>TPAR_L1D1A_AV_dout_nent,
--        nent1=>TPAR_L1D1B_AV_dout_nent,
--        nent2=>TPAR_L1D1C_AV_dout_nent,
--        nent3=>TPAR_L1D1D_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1D1A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L1D1B_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_L1D1C_V_readaddr,
--        addr_arr(39 downto 30)=>TPAR_L1D1D_V_readaddr
--      );

    TPAR_L1D1A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1A_wea_delay,
        addra     => TPAR_L1D1A_writeaddr_delay,
        dina      => TPAR_L1D1A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1A_V_readaddr,
        doutb     => TPAR_L1D1A_V_dout,
        sync_nent => TPAR_L1D1A_start,
        nent_o    => TPAR_L1D1A_AV_dout_nent
      );

    TPAR_L1D1A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1A_wea,
        addra     => TPAR_L1D1A_writeaddr,
        dina      => TPAR_L1D1A_din,
        wea_out       => TPAR_L1D1A_wea_delay,
        addra_out     => TPAR_L1D1A_writeaddr_delay,
        dina_out      => TPAR_L1D1A_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1A_start
      );

    TPAR_L1D1B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1B_wea_delay,
        addra     => TPAR_L1D1B_writeaddr_delay,
        dina      => TPAR_L1D1B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1B_V_readaddr,
        doutb     => TPAR_L1D1B_V_dout,
        sync_nent => TPAR_L1D1B_start,
        nent_o    => TPAR_L1D1B_AV_dout_nent
      );

    TPAR_L1D1B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1B_wea,
        addra     => TPAR_L1D1B_writeaddr,
        dina      => TPAR_L1D1B_din,
        wea_out       => TPAR_L1D1B_wea_delay,
        addra_out     => TPAR_L1D1B_writeaddr_delay,
        dina_out      => TPAR_L1D1B_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1B_start
      );

    TPAR_L1D1C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1C_wea_delay,
        addra     => TPAR_L1D1C_writeaddr_delay,
        dina      => TPAR_L1D1C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1C_V_readaddr,
        doutb     => TPAR_L1D1C_V_dout,
        sync_nent => TPAR_L1D1C_start,
        nent_o    => TPAR_L1D1C_AV_dout_nent
      );

    TPAR_L1D1C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1C_wea,
        addra     => TPAR_L1D1C_writeaddr,
        dina      => TPAR_L1D1C_din,
        wea_out       => TPAR_L1D1C_wea_delay,
        addra_out     => TPAR_L1D1C_writeaddr_delay,
        dina_out      => TPAR_L1D1C_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1C_start
      );

    TPAR_L1D1D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1D_wea_delay,
        addra     => TPAR_L1D1D_writeaddr_delay,
        dina      => TPAR_L1D1D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1D_V_readaddr,
        doutb     => TPAR_L1D1D_V_dout,
        sync_nent => TPAR_L1D1D_start,
        nent_o    => TPAR_L1D1D_AV_dout_nent
      );

    TPAR_L1D1D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1D_wea,
        addra     => TPAR_L1D1D_writeaddr,
        dina      => TPAR_L1D1D_din,
        wea_out       => TPAR_L1D1D_wea_delay,
        addra_out     => TPAR_L1D1D_writeaddr_delay,
        dina_out      => TPAR_L1D1D_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1D_start
      );

    TPARL1D1EFGH_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL1D1EFGH_bx,
        bx_vld => TPARL1D1EFGH_bx_vld
      );

--    MERGE_STREAM_TPARL1D1EFGH : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 4,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL1D1EFGH_bx,
--        bx_in_vld => TPARL1D1EFGH_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L1D1EFGH_stream_V_dout,
--        din0=>TPAR_L1D1E_V_dout,
--        din1=>TPAR_L1D1F_V_dout,
--        din2=>TPAR_L1D1G_V_dout,
--        din3=>TPAR_L1D1H_V_dout,
--        nent0=>TPAR_L1D1E_AV_dout_nent,
--        nent1=>TPAR_L1D1F_AV_dout_nent,
--        nent2=>TPAR_L1D1G_AV_dout_nent,
--        nent3=>TPAR_L1D1H_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L1D1E_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L1D1F_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_L1D1G_V_readaddr,
--        addr_arr(39 downto 30)=>TPAR_L1D1H_V_readaddr
--      );

    TPAR_L1D1E : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1E",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1E_wea_delay,
        addra     => TPAR_L1D1E_writeaddr_delay,
        dina      => TPAR_L1D1E_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1E_V_readaddr,
        doutb     => TPAR_L1D1E_V_dout,
        sync_nent => TPAR_L1D1E_start,
        nent_o    => TPAR_L1D1E_AV_dout_nent
      );

    TPAR_L1D1E_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1E_wea,
        addra     => TPAR_L1D1E_writeaddr,
        dina      => TPAR_L1D1E_din,
        wea_out       => TPAR_L1D1E_wea_delay,
        addra_out     => TPAR_L1D1E_writeaddr_delay,
        dina_out      => TPAR_L1D1E_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1E_start
      );

    TPAR_L1D1F : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1F",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1F_wea_delay,
        addra     => TPAR_L1D1F_writeaddr_delay,
        dina      => TPAR_L1D1F_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1F_V_readaddr,
        doutb     => TPAR_L1D1F_V_dout,
        sync_nent => TPAR_L1D1F_start,
        nent_o    => TPAR_L1D1F_AV_dout_nent
      );

    TPAR_L1D1F_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1F_wea,
        addra     => TPAR_L1D1F_writeaddr,
        dina      => TPAR_L1D1F_din,
        wea_out       => TPAR_L1D1F_wea_delay,
        addra_out     => TPAR_L1D1F_writeaddr_delay,
        dina_out      => TPAR_L1D1F_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1F_start
      );

    TPAR_L1D1G : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1G",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1G_wea_delay,
        addra     => TPAR_L1D1G_writeaddr_delay,
        dina      => TPAR_L1D1G_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1G_V_readaddr,
        doutb     => TPAR_L1D1G_V_dout,
        sync_nent => TPAR_L1D1G_start,
        nent_o    => TPAR_L1D1G_AV_dout_nent
      );

    TPAR_L1D1G_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1G_wea,
        addra     => TPAR_L1D1G_writeaddr,
        dina      => TPAR_L1D1G_din,
        wea_out       => TPAR_L1D1G_wea_delay,
        addra_out     => TPAR_L1D1G_writeaddr_delay,
        dina_out      => TPAR_L1D1G_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1G_start
      );

    TPAR_L1D1H : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L1D1H",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L1D1H_wea_delay,
        addra     => TPAR_L1D1H_writeaddr_delay,
        dina      => TPAR_L1D1H_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L1D1H_V_readaddr,
        doutb     => TPAR_L1D1H_V_dout,
        sync_nent => TPAR_L1D1H_start,
        nent_o    => TPAR_L1D1H_AV_dout_nent
      );

    TPAR_L1D1H_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L1D1H_wea,
        addra     => TPAR_L1D1H_writeaddr,
        dina      => TPAR_L1D1H_din,
        wea_out       => TPAR_L1D1H_wea_delay,
        addra_out     => TPAR_L1D1H_writeaddr_delay,
        dina_out      => TPAR_L1D1H_din_delay,
        done       => TP_done,
        start      => TPAR_L1D1H_start
      );

    TPARL2D1ABCD_STREAM_DELAY : entity work.tf_pipeline_slr_xing
      port map (
        clk => clk,
        bx_out => TP_bx_out,
        bx_out_vld => TP_bx_out_vld,
        bx => TPARL2D1ABCD_bx,
        bx_vld => TPARL2D1ABCD_bx_vld
      );

--    MERGE_STREAM_TPARL2D1ABCD : entity work.tf_merge_streamer
--      generic map (
--        RAM_WIDTH => 73,
--        NUM_PAGES => 8,
--        NUM_INPUTS => 4,
--        NUM_EXTRA_BITS => 2
--      )
--      port map (
--        bx_in => TPARL2D1ABCD_bx,
--        bx_in_vld => TPARL2D1ABCD_bx_vld,
--        rst => '0',
--        clk => clk,
--        merged_dout => MPAR_L2D1ABCD_stream_V_dout,
--        din0=>TPAR_L2D1A_V_dout,
--        din1=>TPAR_L2D1B_V_dout,
--        din2=>TPAR_L2D1C_V_dout,
--        din3=>TPAR_L2D1D_V_dout,
--        nent0=>TPAR_L2D1A_AV_dout_nent,
--        nent1=>TPAR_L2D1B_AV_dout_nent,
--        nent2=>TPAR_L2D1C_AV_dout_nent,
--        nent3=>TPAR_L2D1D_AV_dout_nent,
--        addr_arr(9 downto 0)=>TPAR_L2D1A_V_readaddr,
--        addr_arr(19 downto 10)=>TPAR_L2D1B_V_readaddr,
--        addr_arr(29 downto 20)=>TPAR_L2D1C_V_readaddr,
--        addr_arr(39 downto 30)=>TPAR_L2D1D_V_readaddr
--      );

    TPAR_L2D1A : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2D1A",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2D1A_wea_delay,
        addra     => TPAR_L2D1A_writeaddr_delay,
        dina      => TPAR_L2D1A_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2D1A_V_readaddr,
        doutb     => TPAR_L2D1A_V_dout,
        sync_nent => TPAR_L2D1A_start,
        nent_o    => TPAR_L2D1A_AV_dout_nent
      );

    TPAR_L2D1A_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2D1A_wea,
        addra     => TPAR_L2D1A_writeaddr,
        dina      => TPAR_L2D1A_din,
        wea_out       => TPAR_L2D1A_wea_delay,
        addra_out     => TPAR_L2D1A_writeaddr_delay,
        dina_out      => TPAR_L2D1A_din_delay,
        done       => TP_done,
        start      => TPAR_L2D1A_start
      );

    TPAR_L2D1B : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2D1B",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2D1B_wea_delay,
        addra     => TPAR_L2D1B_writeaddr_delay,
        dina      => TPAR_L2D1B_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2D1B_V_readaddr,
        doutb     => TPAR_L2D1B_V_dout,
        sync_nent => TPAR_L2D1B_start,
        nent_o    => TPAR_L2D1B_AV_dout_nent
      );

    TPAR_L2D1B_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2D1B_wea,
        addra     => TPAR_L2D1B_writeaddr,
        dina      => TPAR_L2D1B_din,
        wea_out       => TPAR_L2D1B_wea_delay,
        addra_out     => TPAR_L2D1B_writeaddr_delay,
        dina_out      => TPAR_L2D1B_din_delay,
        done       => TP_done,
        start      => TPAR_L2D1B_start
      );

    TPAR_L2D1C : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2D1C",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2D1C_wea_delay,
        addra     => TPAR_L2D1C_writeaddr_delay,
        dina      => TPAR_L2D1C_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2D1C_V_readaddr,
        doutb     => TPAR_L2D1C_V_dout,
        sync_nent => TPAR_L2D1C_start,
        nent_o    => TPAR_L2D1C_AV_dout_nent
      );

    TPAR_L2D1C_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2D1C_wea,
        addra     => TPAR_L2D1C_writeaddr,
        dina      => TPAR_L2D1C_din,
        wea_out       => TPAR_L2D1C_wea_delay,
        addra_out     => TPAR_L2D1C_writeaddr_delay,
        dina_out      => TPAR_L2D1C_din_delay,
        done       => TP_done,
        start      => TPAR_L2D1C_start
      );

    TPAR_L2D1D : entity work.tf_mem
      generic map (
        RAM_WIDTH       => 73,
        NUM_PAGES       => 8,
        INIT_FILE       => "",
        INIT_HEX        => true,
        RAM_PERFORMANCE => "HIGH_PERFORMANCE",
        NAME            => "TPAR_L2D1D",
        MEM_TYPE        => "ultra",
        OUT_PIPE_DEPTH  => 2
      )
      port map (
        clka      => clk,
        wea       => TPAR_L2D1D_wea_delay,
        addra     => TPAR_L2D1D_writeaddr_delay,
        dina      => TPAR_L2D1D_din_delay,
        clkb      => clk,
        rstb      => '0',
        regceb    => '1',
        enb       => '1',
        addrb     => TPAR_L2D1D_V_readaddr,
        doutb     => TPAR_L2D1D_V_dout,
        sync_nent => TPAR_L2D1D_start,
        nent_o    => TPAR_L2D1D_AV_dout_nent
      );

    TPAR_L2D1D_DELAY : entity work.tf_pipeline_slr_xing
      generic map (
        NUM_PAGES       => 8,
        RAM_WIDTH       => 73
      )
      port map (
        clk      => clk,
        wea       => TPAR_L2D1D_wea,
        addra     => TPAR_L2D1D_writeaddr,
        dina      => TPAR_L2D1D_din,
        wea_out       => TPAR_L2D1D_wea_delay,
        addra_out     => TPAR_L2D1D_writeaddr_delay,
        dina_out      => TPAR_L2D1D_din_delay,
        done       => TP_done,
        start      => TPAR_L2D1D_start
      );

  LATCH_IR_PS10G_1_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_1_A_bx,
      start => IR_PS10G_1_A_start
  );

  IR_PS10G_1_A : entity work.IR_PS10G_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_1_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => IR_done,
      bx_V          => IR_PS10G_1_A_bx,
      bx_o_V        => IR_bx_out,
      bx_o_V_ap_vld => open,
      hInputStubs_V_dout     => DL_PS10G_1_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_1_A_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_1_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHIA_PS10G_1_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHIA_PS10G_1_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHIA_PS10G_1_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIB_PS10G_1_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIB_PS10G_1_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIB_PS10G_1_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L1PHIC_PS10G_1_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L1PHIC_PS10G_1_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L1PHIC_PS10G_1_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L1PHID_PS10G_1_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L1PHID_PS10G_1_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L1PHID_PS10G_1_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_L1PHIE_PS10G_1_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_L1PHIE_PS10G_1_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_L1PHIE_PS10G_1_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D1PHIA_PS10G_1_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D1PHIA_PS10G_1_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D1PHIA_PS10G_1_A_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D1PHIB_PS10G_1_A_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D1PHIB_PS10G_1_A_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D1PHIB_PS10G_1_A_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D1PHIC_PS10G_1_A_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D1PHIC_PS10G_1_A_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D1PHIC_PS10G_1_A_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D3PHIA_PS10G_1_A_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D3PHIA_PS10G_1_A_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D3PHIA_PS10G_1_A_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D3PHIB_PS10G_1_A_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D3PHIB_PS10G_1_A_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D3PHIB_PS10G_1_A_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D3PHIC_PS10G_1_A_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D3PHIC_PS10G_1_A_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D3PHIC_PS10G_1_A_din,
      hOutputStubs_11_dataarray_data_V_ce0       => open,
      hOutputStubs_11_dataarray_data_V_we0       => IL_D5PHIA_PS10G_1_A_wea,
      hOutputStubs_11_dataarray_data_V_address0  => IL_D5PHIA_PS10G_1_A_writeaddr,
      hOutputStubs_11_dataarray_data_V_d0        => IL_D5PHIA_PS10G_1_A_din,
      hOutputStubs_12_dataarray_data_V_ce0       => open,
      hOutputStubs_12_dataarray_data_V_we0       => IL_D5PHIB_PS10G_1_A_wea,
      hOutputStubs_12_dataarray_data_V_address0  => IL_D5PHIB_PS10G_1_A_writeaddr,
      hOutputStubs_12_dataarray_data_V_d0        => IL_D5PHIB_PS10G_1_A_din,
      hOutputStubs_13_dataarray_data_V_ce0       => open,
      hOutputStubs_13_dataarray_data_V_we0       => IL_D5PHIC_PS10G_1_A_wea,
      hOutputStubs_13_dataarray_data_V_address0  => IL_D5PHIC_PS10G_1_A_writeaddr,
      hOutputStubs_13_dataarray_data_V_d0        => IL_D5PHIC_PS10G_1_A_din,
      hLinkWord_V => "10001010011000100011",
      hPhBnWord_V => "00000111000001110000011100011111"
  );

  LATCH_IR_PS10G_1_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_1_B_bx,
      start => IR_PS10G_1_B_start
  );

  IR_PS10G_1_B : entity work.IR_PS10G_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_1_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS10G_1_B_bx,
      hInputStubs_V_dout     => DL_PS10G_1_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_1_B_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_1_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHIG_PS10G_1_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHIG_PS10G_1_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHIG_PS10G_1_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIH_PS10G_1_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIH_PS10G_1_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIH_PS10G_1_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHIB_PS10G_1_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHIB_PS10G_1_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHIB_PS10G_1_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D1PHIC_PS10G_1_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D1PHIC_PS10G_1_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D1PHIC_PS10G_1_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D1PHID_PS10G_1_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D1PHID_PS10G_1_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D1PHID_PS10G_1_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHIB_PS10G_1_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHIB_PS10G_1_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHIB_PS10G_1_B_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D3PHIC_PS10G_1_B_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D3PHIC_PS10G_1_B_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D3PHIC_PS10G_1_B_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D3PHID_PS10G_1_B_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D3PHID_PS10G_1_B_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D3PHID_PS10G_1_B_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D5PHIB_PS10G_1_B_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D5PHIB_PS10G_1_B_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D5PHIB_PS10G_1_B_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D5PHIC_PS10G_1_B_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D5PHIC_PS10G_1_B_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D5PHIC_PS10G_1_B_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D5PHID_PS10G_1_B_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D5PHID_PS10G_1_B_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D5PHID_PS10G_1_B_din,
      hLinkWord_V => "10001010011000100011",
      hPhBnWord_V => "00001110000011100000111011000000"
  );

  LATCH_IR_PS10G_2_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_2_A_bx,
      start => IR_PS10G_2_A_start
  );

  IR_PS10G_2_A : entity work.IR_PS10G_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_2_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS10G_2_A_bx,
      hInputStubs_V_dout     => DL_PS10G_2_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_2_A_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_2_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHIA_PS10G_2_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHIA_PS10G_2_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHIA_PS10G_2_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIB_PS10G_2_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIB_PS10G_2_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIB_PS10G_2_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L1PHIC_PS10G_2_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L1PHIC_PS10G_2_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L1PHIC_PS10G_2_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L1PHID_PS10G_2_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L1PHID_PS10G_2_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L1PHID_PS10G_2_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_L1PHIE_PS10G_2_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_L1PHIE_PS10G_2_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_L1PHIE_PS10G_2_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHIA_PS10G_2_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHIA_PS10G_2_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHIA_PS10G_2_A_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D2PHIB_PS10G_2_A_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D2PHIB_PS10G_2_A_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D2PHIB_PS10G_2_A_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D2PHIC_PS10G_2_A_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D2PHIC_PS10G_2_A_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D2PHIC_PS10G_2_A_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D4PHIA_PS10G_2_A_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D4PHIA_PS10G_2_A_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D4PHIA_PS10G_2_A_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D4PHIB_PS10G_2_A_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D4PHIB_PS10G_2_A_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D4PHIB_PS10G_2_A_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D4PHIC_PS10G_2_A_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D4PHIC_PS10G_2_A_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D4PHIC_PS10G_2_A_din,
      hLinkWord_V => "01100000100001000011",
      hPhBnWord_V => "00000000000001110000011100011111"
  );

  LATCH_IR_PS10G_2_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_2_B_bx,
      start => IR_PS10G_2_B_start
  );

  IR_PS10G_2_B : entity work.IR_PS10G_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_2_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS10G_2_B_bx,
      hInputStubs_V_dout     => DL_PS10G_2_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_2_B_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_2_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHID_PS10G_2_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHID_PS10G_2_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHID_PS10G_2_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIE_PS10G_2_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIE_PS10G_2_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIE_PS10G_2_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L1PHIF_PS10G_2_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L1PHIF_PS10G_2_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L1PHIF_PS10G_2_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L1PHIG_PS10G_2_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L1PHIG_PS10G_2_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L1PHIG_PS10G_2_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_L1PHIH_PS10G_2_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_L1PHIH_PS10G_2_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_L1PHIH_PS10G_2_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHIB_PS10G_2_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHIB_PS10G_2_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHIB_PS10G_2_B_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D2PHIC_PS10G_2_B_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D2PHIC_PS10G_2_B_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D2PHIC_PS10G_2_B_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D2PHID_PS10G_2_B_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D2PHID_PS10G_2_B_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D2PHID_PS10G_2_B_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D4PHIB_PS10G_2_B_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D4PHIB_PS10G_2_B_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D4PHIB_PS10G_2_B_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D4PHIC_PS10G_2_B_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D4PHIC_PS10G_2_B_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D4PHIC_PS10G_2_B_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D4PHID_PS10G_2_B_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D4PHID_PS10G_2_B_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D4PHID_PS10G_2_B_din,
      hLinkWord_V => "01100000100001000011",
      hPhBnWord_V => "00000000000011100000111011111000"
  );

  LATCH_IR_PS10G_3_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_3_A_bx,
      start => IR_PS10G_3_A_start
  );

  IR_PS10G_3_A : entity work.IR_PS10G_3_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_3_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS10G_3_A_bx,
      hInputStubs_V_dout     => DL_PS10G_3_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_3_A_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_3_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L2PHIA_PS10G_3_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L2PHIA_PS10G_3_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L2PHIA_PS10G_3_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L2PHIB_PS10G_3_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L2PHIB_PS10G_3_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L2PHIB_PS10G_3_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L2PHIC_PS10G_3_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L2PHIC_PS10G_3_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L2PHIC_PS10G_3_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIA_PS10G_3_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIA_PS10G_3_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIA_PS10G_3_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHIB_PS10G_3_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHIB_PS10G_3_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHIB_PS10G_3_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHIC_PS10G_3_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHIC_PS10G_3_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHIC_PS10G_3_A_din,
      hLinkWord_V => "01000000000001000101",
      hPhBnWord_V => "00000000000000000000011100000111"
  );

  LATCH_IR_PS10G_3_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_3_B_bx,
      start => IR_PS10G_3_B_start
  );

  IR_PS10G_3_B : entity work.IR_PS10G_3_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_3_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS10G_3_B_bx,
      hInputStubs_V_dout     => DL_PS10G_3_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_3_B_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_3_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L2PHIB_PS10G_3_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L2PHIB_PS10G_3_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L2PHIB_PS10G_3_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L2PHIC_PS10G_3_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L2PHIC_PS10G_3_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L2PHIC_PS10G_3_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L2PHID_PS10G_3_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L2PHID_PS10G_3_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L2PHID_PS10G_3_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIB_PS10G_3_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIB_PS10G_3_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIB_PS10G_3_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHIC_PS10G_3_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHIC_PS10G_3_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHIC_PS10G_3_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHID_PS10G_3_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHID_PS10G_3_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHID_PS10G_3_B_din,
      hLinkWord_V => "01000000000001000101",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_PS10G_4_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_4_A_bx,
      start => IR_PS10G_4_A_start
  );

  IR_PS10G_4_A : entity work.IR_PS10G_4_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_4_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS10G_4_A_bx,
      hInputStubs_V_dout     => DL_PS10G_4_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_4_A_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_4_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIA_PS10G_4_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIA_PS10G_4_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIA_PS10G_4_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIB_PS10G_4_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIB_PS10G_4_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIB_PS10G_4_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHIC_PS10G_4_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHIC_PS10G_4_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHIC_PS10G_4_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIA_PS10G_4_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIA_PS10G_4_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIA_PS10G_4_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIB_PS10G_4_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIB_PS10G_4_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIB_PS10G_4_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHIC_PS10G_4_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHIC_PS10G_4_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHIC_PS10G_4_A_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D5PHIA_PS10G_4_A_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D5PHIA_PS10G_4_A_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D5PHIA_PS10G_4_A_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D5PHIB_PS10G_4_A_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D5PHIB_PS10G_4_A_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D5PHIB_PS10G_4_A_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D5PHIC_PS10G_4_A_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D5PHIC_PS10G_4_A_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D5PHIC_PS10G_4_A_din,
      hLinkWord_V => "01100000101001100010",
      hPhBnWord_V => "00000000000001110000011100000111"
  );

  LATCH_IR_PS10G_4_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS10G_4_B_bx,
      start => IR_PS10G_4_B_start
  );

  IR_PS10G_4_B : entity work.IR_PS10G_4_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS10G_4_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS10G_4_B_bx,
      hInputStubs_V_dout     => DL_PS10G_4_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS10G_4_B_link_empty_neg,
      hInputStubs_V_read     => DL_PS10G_4_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIB_PS10G_4_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIB_PS10G_4_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIB_PS10G_4_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIC_PS10G_4_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIC_PS10G_4_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIC_PS10G_4_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHID_PS10G_4_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHID_PS10G_4_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHID_PS10G_4_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIB_PS10G_4_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIB_PS10G_4_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIB_PS10G_4_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIC_PS10G_4_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIC_PS10G_4_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIC_PS10G_4_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHID_PS10G_4_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHID_PS10G_4_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHID_PS10G_4_B_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D5PHIB_PS10G_4_B_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D5PHIB_PS10G_4_B_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D5PHIB_PS10G_4_B_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D5PHIC_PS10G_4_B_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D5PHIC_PS10G_4_B_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D5PHIC_PS10G_4_B_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D5PHID_PS10G_4_B_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D5PHID_PS10G_4_B_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D5PHID_PS10G_4_B_din,
      hLinkWord_V => "01100000101001100010",
      hPhBnWord_V => "00000000000011100000111000001110"
  );

  LATCH_IR_PS_1_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS_1_A_bx,
      start => IR_PS_1_A_start
  );

  IR_PS_1_A : entity work.IR_PS_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS_1_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS_1_A_bx,
      hInputStubs_V_dout     => DL_PS_1_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS_1_A_link_empty_neg,
      hInputStubs_V_read     => DL_PS_1_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIA_PS_1_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIA_PS_1_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIA_PS_1_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHIB_PS_1_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHIB_PS_1_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHIB_PS_1_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D2PHIA_PS_1_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D2PHIA_PS_1_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D2PHIA_PS_1_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIB_PS_1_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIB_PS_1_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIB_PS_1_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHIC_PS_1_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHIC_PS_1_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHIC_PS_1_A_din,
      hLinkWord_V => "01000000000001000111",
      hPhBnWord_V => "00000000000000000000011100000011"
  );

  LATCH_IR_PS_1_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS_1_B_bx,
      start => IR_PS_1_B_start
  );

  IR_PS_1_B : entity work.IR_PS_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS_1_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS_1_B_bx,
      hInputStubs_V_dout     => DL_PS_1_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS_1_B_link_empty_neg,
      hInputStubs_V_read     => DL_PS_1_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIC_PS_1_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIC_PS_1_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIC_PS_1_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHID_PS_1_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHID_PS_1_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHID_PS_1_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D2PHIB_PS_1_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D2PHIB_PS_1_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D2PHIB_PS_1_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIC_PS_1_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIC_PS_1_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIC_PS_1_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHID_PS_1_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHID_PS_1_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHID_PS_1_B_din,
      hLinkWord_V => "01000000000001000111",
      hPhBnWord_V => "00000000000000000000111000001100"
  );

  LATCH_IR_PS_2_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS_2_A_bx,
      start => IR_PS_2_A_start
  );

  IR_PS_2_A : entity work.IR_PS_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS_2_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS_2_A_bx,
      hInputStubs_V_dout     => DL_PS_2_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS_2_A_link_empty_neg,
      hInputStubs_V_read     => DL_PS_2_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIA_PS_2_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIA_PS_2_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIA_PS_2_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHIB_PS_2_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHIB_PS_2_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHIB_PS_2_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D4PHIA_PS_2_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D4PHIA_PS_2_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D4PHIA_PS_2_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIB_PS_2_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIB_PS_2_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIB_PS_2_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIC_PS_2_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIC_PS_2_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIC_PS_2_A_din,
      hLinkWord_V => "01000000000010000111",
      hPhBnWord_V => "00000000000000000000011100000011"
  );

  LATCH_IR_PS_2_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_PS_2_B_bx,
      start => IR_PS_2_B_start
  );

  IR_PS_2_B : entity work.IR_PS_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_PS_2_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_PS_2_B_bx,
      hInputStubs_V_dout     => DL_PS_2_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_PS_2_B_link_empty_neg,
      hInputStubs_V_read     => DL_PS_2_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIB_PS_2_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIB_PS_2_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIB_PS_2_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHIC_PS_2_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHIC_PS_2_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHIC_PS_2_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L3PHID_PS_2_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L3PHID_PS_2_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L3PHID_PS_2_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIB_PS_2_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIB_PS_2_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIB_PS_2_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIC_PS_2_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIC_PS_2_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIC_PS_2_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D4PHID_PS_2_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D4PHID_PS_2_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D4PHID_PS_2_B_din,
      hLinkWord_V => "01000000000010000111",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_negPS10G_1_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_1_A_bx,
      start => IR_negPS10G_1_A_start
  );

  IR_negPS10G_1_A : entity work.IR_negPS10G_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_1_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_1_A_bx,
      hInputStubs_V_dout     => DL_negPS10G_1_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_1_A_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_1_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHIA_negPS10G_1_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHIA_negPS10G_1_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHIA_negPS10G_1_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIB_negPS10G_1_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIB_negPS10G_1_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIB_negPS10G_1_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHIA_negPS10G_1_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHIA_negPS10G_1_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHIA_negPS10G_1_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D1PHIB_negPS10G_1_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_1_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D1PHIB_negPS10G_1_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D1PHIC_negPS10G_1_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_1_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D1PHIC_negPS10G_1_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHIA_negPS10G_1_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHIA_negPS10G_1_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHIA_negPS10G_1_A_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D3PHIB_negPS10G_1_A_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_1_A_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D3PHIB_negPS10G_1_A_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D3PHIC_negPS10G_1_A_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_1_A_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D3PHIC_negPS10G_1_A_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D5PHIA_negPS10G_1_A_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D5PHIA_negPS10G_1_A_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D5PHIA_negPS10G_1_A_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D5PHIB_negPS10G_1_A_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_1_A_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D5PHIB_negPS10G_1_A_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D5PHIC_negPS10G_1_A_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_1_A_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D5PHIC_negPS10G_1_A_din,
      hLinkWord_V => "10001010011000100011",
      hPhBnWord_V => "00000111000001110000011100000011"
  );

  LATCH_IR_negPS10G_1_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_1_B_bx,
      start => IR_negPS10G_1_B_start
  );

  IR_negPS10G_1_B : entity work.IR_negPS10G_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_1_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_1_B_bx,
      hInputStubs_V_dout     => DL_negPS10G_1_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_1_B_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_1_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHID_negPS10G_1_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHID_negPS10G_1_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHID_negPS10G_1_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIE_negPS10G_1_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIE_negPS10G_1_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIE_negPS10G_1_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L1PHIF_negPS10G_1_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L1PHIF_negPS10G_1_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L1PHIF_negPS10G_1_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L1PHIG_negPS10G_1_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L1PHIG_negPS10G_1_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L1PHIG_negPS10G_1_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D1PHIB_negPS10G_1_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_1_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D1PHIB_negPS10G_1_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D1PHIC_negPS10G_1_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_1_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D1PHIC_negPS10G_1_B_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D1PHID_negPS10G_1_B_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D1PHID_negPS10G_1_B_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D1PHID_negPS10G_1_B_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D3PHIB_negPS10G_1_B_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_1_B_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D3PHIB_negPS10G_1_B_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D3PHIC_negPS10G_1_B_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_1_B_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D3PHIC_negPS10G_1_B_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D3PHID_negPS10G_1_B_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D3PHID_negPS10G_1_B_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D3PHID_negPS10G_1_B_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D5PHIB_negPS10G_1_B_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_1_B_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D5PHIB_negPS10G_1_B_din,
      hOutputStubs_11_dataarray_data_V_ce0       => open,
      hOutputStubs_11_dataarray_data_V_we0       => IL_D5PHIC_negPS10G_1_B_wea,
      hOutputStubs_11_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_1_B_writeaddr,
      hOutputStubs_11_dataarray_data_V_d0        => IL_D5PHIC_negPS10G_1_B_din,
      hOutputStubs_12_dataarray_data_V_ce0       => open,
      hOutputStubs_12_dataarray_data_V_we0       => IL_D5PHID_negPS10G_1_B_wea,
      hOutputStubs_12_dataarray_data_V_address0  => IL_D5PHID_negPS10G_1_B_writeaddr,
      hOutputStubs_12_dataarray_data_V_d0        => IL_D5PHID_negPS10G_1_B_din,
      hLinkWord_V => "10001010011000100011",
      hPhBnWord_V => "00001110000011100000111001111000"
  );

  LATCH_IR_negPS10G_2_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_2_A_bx,
      start => IR_negPS10G_2_A_start
  );

  IR_negPS10G_2_A : entity work.IR_negPS10G_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_2_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_2_A_bx,
      hInputStubs_V_dout     => DL_negPS10G_2_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_2_A_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_2_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHIA_negPS10G_2_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHIA_negPS10G_2_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHIA_negPS10G_2_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIB_negPS10G_2_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIB_negPS10G_2_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIB_negPS10G_2_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L1PHIC_negPS10G_2_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L1PHIC_negPS10G_2_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L1PHIC_negPS10G_2_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L1PHID_negPS10G_2_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L1PHID_negPS10G_2_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L1PHID_negPS10G_2_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_L1PHIE_negPS10G_2_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_L1PHIE_negPS10G_2_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_L1PHIE_negPS10G_2_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHIA_negPS10G_2_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHIA_negPS10G_2_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHIA_negPS10G_2_A_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D2PHIB_negPS10G_2_A_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_2_A_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D2PHIB_negPS10G_2_A_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D2PHIC_negPS10G_2_A_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_2_A_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D2PHIC_negPS10G_2_A_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D4PHIA_negPS10G_2_A_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D4PHIA_negPS10G_2_A_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D4PHIA_negPS10G_2_A_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D4PHIB_negPS10G_2_A_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D4PHIB_negPS10G_2_A_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D4PHIB_negPS10G_2_A_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D4PHIC_negPS10G_2_A_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D4PHIC_negPS10G_2_A_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D4PHIC_negPS10G_2_A_din,
      hLinkWord_V => "01100000100001000011",
      hPhBnWord_V => "00000000000001110000011100011111"
  );

  LATCH_IR_negPS10G_2_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_2_B_bx,
      start => IR_negPS10G_2_B_start
  );

  IR_negPS10G_2_B : entity work.IR_negPS10G_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_2_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_2_B_bx,
      hInputStubs_V_dout     => DL_negPS10G_2_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_2_B_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_2_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L1PHID_negPS10G_2_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L1PHID_negPS10G_2_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L1PHID_negPS10G_2_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L1PHIE_negPS10G_2_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L1PHIE_negPS10G_2_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L1PHIE_negPS10G_2_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L1PHIF_negPS10G_2_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L1PHIF_negPS10G_2_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L1PHIF_negPS10G_2_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L1PHIG_negPS10G_2_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L1PHIG_negPS10G_2_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L1PHIG_negPS10G_2_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_L1PHIH_negPS10G_2_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_L1PHIH_negPS10G_2_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_L1PHIH_negPS10G_2_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHIB_negPS10G_2_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_2_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHIB_negPS10G_2_B_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D2PHIC_negPS10G_2_B_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_2_B_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D2PHIC_negPS10G_2_B_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D2PHID_negPS10G_2_B_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D2PHID_negPS10G_2_B_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D2PHID_negPS10G_2_B_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D4PHIB_negPS10G_2_B_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D4PHIB_negPS10G_2_B_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D4PHIB_negPS10G_2_B_din,
      hOutputStubs_9_dataarray_data_V_ce0       => open,
      hOutputStubs_9_dataarray_data_V_we0       => IL_D4PHIC_negPS10G_2_B_wea,
      hOutputStubs_9_dataarray_data_V_address0  => IL_D4PHIC_negPS10G_2_B_writeaddr,
      hOutputStubs_9_dataarray_data_V_d0        => IL_D4PHIC_negPS10G_2_B_din,
      hOutputStubs_10_dataarray_data_V_ce0       => open,
      hOutputStubs_10_dataarray_data_V_we0       => IL_D4PHID_negPS10G_2_B_wea,
      hOutputStubs_10_dataarray_data_V_address0  => IL_D4PHID_negPS10G_2_B_writeaddr,
      hOutputStubs_10_dataarray_data_V_d0        => IL_D4PHID_negPS10G_2_B_din,
      hLinkWord_V => "01100000100001000011",
      hPhBnWord_V => "00000000000011100000111011111000"
  );

  LATCH_IR_negPS10G_3_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_3_A_bx,
      start => IR_negPS10G_3_A_start
  );

  IR_negPS10G_3_A : entity work.IR_negPS10G_3_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_3_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_3_A_bx,
      hInputStubs_V_dout     => DL_negPS10G_3_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_3_A_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_3_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L2PHIA_negPS10G_3_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L2PHIA_negPS10G_3_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L2PHIA_negPS10G_3_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L2PHIB_negPS10G_3_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L2PHIB_negPS10G_3_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L2PHIB_negPS10G_3_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L2PHIC_negPS10G_3_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L2PHIC_negPS10G_3_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L2PHIC_negPS10G_3_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIA_negPS10G_3_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIA_negPS10G_3_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIA_negPS10G_3_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHIB_negPS10G_3_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_3_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHIB_negPS10G_3_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHIC_negPS10G_3_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_3_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHIC_negPS10G_3_A_din,
      hLinkWord_V => "01000000000001000101",
      hPhBnWord_V => "00000000000000000000011100000111"
  );

  LATCH_IR_negPS10G_3_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_3_B_bx,
      start => IR_negPS10G_3_B_start
  );

  IR_negPS10G_3_B : entity work.IR_negPS10G_3_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_3_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_3_B_bx,
      hInputStubs_V_dout     => DL_negPS10G_3_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_3_B_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_3_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L2PHIB_negPS10G_3_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L2PHIB_negPS10G_3_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L2PHIB_negPS10G_3_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L2PHIC_negPS10G_3_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L2PHIC_negPS10G_3_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L2PHIC_negPS10G_3_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L2PHID_negPS10G_3_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L2PHID_negPS10G_3_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L2PHID_negPS10G_3_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIB_negPS10G_3_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_3_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIB_negPS10G_3_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHIC_negPS10G_3_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_3_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHIC_negPS10G_3_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHID_negPS10G_3_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHID_negPS10G_3_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHID_negPS10G_3_B_din,
      hLinkWord_V => "01000000000001000101",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_negPS10G_4_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_4_A_bx,
      start => IR_negPS10G_4_A_start
  );

  IR_negPS10G_4_A : entity work.IR_negPS10G_4_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_4_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_4_A_bx,
      hInputStubs_V_dout     => DL_negPS10G_4_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_4_A_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_4_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIA_negPS10G_4_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIA_negPS10G_4_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIA_negPS10G_4_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIB_negPS10G_4_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_4_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIB_negPS10G_4_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHIC_negPS10G_4_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_4_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHIC_negPS10G_4_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIA_negPS10G_4_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIA_negPS10G_4_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIA_negPS10G_4_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIB_negPS10G_4_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_4_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIB_negPS10G_4_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHIC_negPS10G_4_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_4_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHIC_negPS10G_4_A_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D5PHIA_negPS10G_4_A_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D5PHIA_negPS10G_4_A_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D5PHIA_negPS10G_4_A_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D5PHIB_negPS10G_4_A_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_4_A_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D5PHIB_negPS10G_4_A_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D5PHIC_negPS10G_4_A_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_4_A_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D5PHIC_negPS10G_4_A_din,
      hLinkWord_V => "01100000101001100010",
      hPhBnWord_V => "00000000000001110000011100000111"
  );

  LATCH_IR_negPS10G_4_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS10G_4_B_bx,
      start => IR_negPS10G_4_B_start
  );

  IR_negPS10G_4_B : entity work.IR_negPS10G_4_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS10G_4_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS10G_4_B_bx,
      hInputStubs_V_dout     => DL_negPS10G_4_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS10G_4_B_link_empty_neg,
      hInputStubs_V_read     => DL_negPS10G_4_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIB_negPS10G_4_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_4_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIB_negPS10G_4_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIC_negPS10G_4_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_4_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIC_negPS10G_4_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHID_negPS10G_4_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHID_negPS10G_4_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHID_negPS10G_4_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIB_negPS10G_4_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_4_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIB_negPS10G_4_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIC_negPS10G_4_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_4_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIC_negPS10G_4_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHID_negPS10G_4_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHID_negPS10G_4_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHID_negPS10G_4_B_din,
      hOutputStubs_6_dataarray_data_V_ce0       => open,
      hOutputStubs_6_dataarray_data_V_we0       => IL_D5PHIB_negPS10G_4_B_wea,
      hOutputStubs_6_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_4_B_writeaddr,
      hOutputStubs_6_dataarray_data_V_d0        => IL_D5PHIB_negPS10G_4_B_din,
      hOutputStubs_7_dataarray_data_V_ce0       => open,
      hOutputStubs_7_dataarray_data_V_we0       => IL_D5PHIC_negPS10G_4_B_wea,
      hOutputStubs_7_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_4_B_writeaddr,
      hOutputStubs_7_dataarray_data_V_d0        => IL_D5PHIC_negPS10G_4_B_din,
      hOutputStubs_8_dataarray_data_V_ce0       => open,
      hOutputStubs_8_dataarray_data_V_we0       => IL_D5PHID_negPS10G_4_B_wea,
      hOutputStubs_8_dataarray_data_V_address0  => IL_D5PHID_negPS10G_4_B_writeaddr,
      hOutputStubs_8_dataarray_data_V_d0        => IL_D5PHID_negPS10G_4_B_din,
      hLinkWord_V => "01100000101001100010",
      hPhBnWord_V => "00000000000011100000111000001110"
  );

  LATCH_IR_negPS_1_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS_1_A_bx,
      start => IR_negPS_1_A_start
  );

  IR_negPS_1_A : entity work.IR_negPS_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS_1_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS_1_A_bx,
      hInputStubs_V_dout     => DL_negPS_1_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS_1_A_link_empty_neg,
      hInputStubs_V_read     => DL_negPS_1_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIA_negPS_1_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIA_negPS_1_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIA_negPS_1_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHIB_negPS_1_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHIB_negPS_1_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHIB_negPS_1_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D2PHIA_negPS_1_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D2PHIA_negPS_1_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D2PHIA_negPS_1_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIB_negPS_1_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIB_negPS_1_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIB_negPS_1_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHIC_negPS_1_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHIC_negPS_1_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHIC_negPS_1_A_din,
      hLinkWord_V => "01000000000001000111",
      hPhBnWord_V => "00000000000000000000011100000011"
  );

  LATCH_IR_negPS_1_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS_1_B_bx,
      start => IR_negPS_1_B_start
  );

  IR_negPS_1_B : entity work.IR_negPS_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS_1_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS_1_B_bx,
      hInputStubs_V_dout     => DL_negPS_1_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS_1_B_link_empty_neg,
      hInputStubs_V_read     => DL_negPS_1_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIB_negPS_1_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIB_negPS_1_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIB_negPS_1_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHIC_negPS_1_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHIC_negPS_1_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHIC_negPS_1_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L3PHID_negPS_1_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L3PHID_negPS_1_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L3PHID_negPS_1_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D2PHIB_negPS_1_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D2PHIB_negPS_1_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D2PHIB_negPS_1_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D2PHIC_negPS_1_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D2PHIC_negPS_1_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D2PHIC_negPS_1_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D2PHID_negPS_1_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D2PHID_negPS_1_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D2PHID_negPS_1_B_din,
      hLinkWord_V => "01000000000001000111",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_negPS_2_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS_2_A_bx,
      start => IR_negPS_2_A_start
  );

  IR_negPS_2_A : entity work.IR_negPS_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS_2_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS_2_A_bx,
      hInputStubs_V_dout     => DL_negPS_2_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS_2_A_link_empty_neg,
      hInputStubs_V_read     => DL_negPS_2_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIA_negPS_2_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIA_negPS_2_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIA_negPS_2_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHIB_negPS_2_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHIB_negPS_2_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHIB_negPS_2_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D4PHIA_negPS_2_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D4PHIA_negPS_2_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D4PHIA_negPS_2_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIB_negPS_2_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIB_negPS_2_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIB_negPS_2_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIC_negPS_2_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIC_negPS_2_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIC_negPS_2_A_din,
      hLinkWord_V => "01000000000010000111",
      hPhBnWord_V => "00000000000000000000011100000011"
  );

  LATCH_IR_negPS_2_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_negPS_2_B_bx,
      start => IR_negPS_2_B_start
  );

  IR_negPS_2_B : entity work.IR_negPS_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_negPS_2_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_negPS_2_B_bx,
      hInputStubs_V_dout     => DL_negPS_2_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_negPS_2_B_link_empty_neg,
      hInputStubs_V_read     => DL_negPS_2_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L3PHIB_negPS_2_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L3PHIB_negPS_2_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L3PHIB_negPS_2_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L3PHIC_negPS_2_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L3PHIC_negPS_2_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L3PHIC_negPS_2_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L3PHID_negPS_2_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L3PHID_negPS_2_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L3PHID_negPS_2_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIB_negPS_2_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIB_negPS_2_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIB_negPS_2_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIC_negPS_2_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIC_negPS_2_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIC_negPS_2_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D4PHID_negPS_2_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D4PHID_negPS_2_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D4PHID_negPS_2_B_din,
      hLinkWord_V => "01000000000010000111",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_2S_1_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_1_A_bx,
      start => IR_2S_1_A_start
  );

  IR_2S_1_A : entity work.IR_2S_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_1_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_1_A_bx,
      hInputStubs_V_dout     => DL_twoS_1_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_1_A_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_1_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L4PHIA_2S_1_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L4PHIA_2S_1_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L4PHIA_2S_1_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L4PHIB_2S_1_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L4PHIB_2S_1_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L4PHIB_2S_1_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L4PHIC_2S_1_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L4PHIC_2S_1_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L4PHIC_2S_1_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L5PHIA_2S_1_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L5PHIA_2S_1_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L5PHIA_2S_1_A_din,
      hLinkWord_V => "01010000000010111001",
      hPhBnWord_V => "00000000000000000000000100000111"
  );

  LATCH_IR_2S_1_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_1_B_bx,
      start => IR_2S_1_B_start
  );

  IR_2S_1_B : entity work.IR_2S_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_1_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_1_B_bx,
      hInputStubs_V_dout     => DL_twoS_1_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_1_B_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_1_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L4PHIB_2S_1_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L4PHIB_2S_1_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L4PHIB_2S_1_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L4PHIC_2S_1_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L4PHIC_2S_1_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L4PHIC_2S_1_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L4PHID_2S_1_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L4PHID_2S_1_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L4PHID_2S_1_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L5PHID_2S_1_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L5PHID_2S_1_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L5PHID_2S_1_B_din,
      hLinkWord_V => "01010000000010111001",
      hPhBnWord_V => "00000000000000000000100000001110"
  );

  LATCH_IR_2S_2_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_2_A_bx,
      start => IR_2S_2_A_start
  );

  IR_2S_2_A : entity work.IR_2S_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_2_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_2_A_bx,
      hInputStubs_V_dout     => DL_twoS_2_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_2_A_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_2_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L5PHIA_2S_2_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L5PHIA_2S_2_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L5PHIA_2S_2_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L5PHIB_2S_2_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L5PHIB_2S_2_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L5PHIB_2S_2_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L5PHIC_2S_2_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L5PHIC_2S_2_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L5PHIC_2S_2_A_din,
      hLinkWord_V => "00110000000000001011",
      hPhBnWord_V => "00000000000000000000000000000111"
  );

  LATCH_IR_2S_2_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_2_B_bx,
      start => IR_2S_2_B_start
  );

  IR_2S_2_B : entity work.IR_2S_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_2_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_2_B_bx,
      hInputStubs_V_dout     => DL_twoS_2_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_2_B_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_2_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L5PHIB_2S_2_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L5PHIB_2S_2_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L5PHIB_2S_2_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L5PHIC_2S_2_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L5PHIC_2S_2_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L5PHIC_2S_2_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L5PHID_2S_2_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L5PHID_2S_2_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L5PHID_2S_2_B_din,
      hLinkWord_V => "00110000000000001011",
      hPhBnWord_V => "00000000000000000000000000001110"
  );

  LATCH_IR_2S_3_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_3_A_bx,
      start => IR_2S_3_A_start
  );

  IR_2S_3_A : entity work.IR_2S_3_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_3_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_3_A_bx,
      hInputStubs_V_dout     => DL_twoS_3_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_3_A_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_3_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIA_2S_3_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIA_2S_3_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIA_2S_3_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHIB_2S_3_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHIB_2S_3_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHIB_2S_3_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L6PHIC_2S_3_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L6PHIC_2S_3_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L6PHIC_2S_3_A_din,
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "00000000000000000000000000000111"
  );

  LATCH_IR_2S_3_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_3_B_bx,
      start => IR_2S_3_B_start
  );

  IR_2S_3_B : entity work.IR_2S_3_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_3_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_3_B_bx,
      hInputStubs_V_dout     => DL_twoS_3_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_3_B_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_3_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIC_2S_3_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIC_2S_3_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIC_2S_3_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHID_2S_3_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHID_2S_3_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHID_2S_3_B_din,
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "00000000000000000000000000001100"
  );

  LATCH_IR_2S_4_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_4_A_bx,
      start => IR_2S_4_A_start
  );

  IR_2S_4_A : entity work.IR_2S_4_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_4_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_4_A_bx,
      hInputStubs_V_dout     => DL_twoS_4_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_4_A_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_4_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIA_2S_4_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIA_2S_4_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIA_2S_4_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHIB_2S_4_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHIB_2S_4_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHIB_2S_4_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D3PHIA_2S_4_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D3PHIA_2S_4_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D3PHIA_2S_4_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIB_2S_4_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIB_2S_4_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIB_2S_4_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIC_2S_4_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIC_2S_4_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIC_2S_4_A_din,
      hLinkWord_V => "01010000000001101101",
      hPhBnWord_V => "00000000000000000000011100000011"
  );

  LATCH_IR_2S_4_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_4_B_bx,
      start => IR_2S_4_B_start
  );

  IR_2S_4_B : entity work.IR_2S_4_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_4_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_4_B_bx,
      hInputStubs_V_dout     => DL_twoS_4_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_4_B_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_4_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIB_2S_4_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIB_2S_4_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIB_2S_4_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHIC_2S_4_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHIC_2S_4_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHIC_2S_4_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L6PHID_2S_4_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L6PHID_2S_4_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L6PHID_2S_4_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIB_2S_4_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIB_2S_4_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIB_2S_4_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIC_2S_4_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIC_2S_4_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIC_2S_4_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHID_2S_4_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHID_2S_4_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHID_2S_4_B_din,
      hLinkWord_V => "01010000000001101101",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_2S_5_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_5_A_bx,
      start => IR_2S_5_A_start
  );

  IR_2S_5_A : entity work.IR_2S_5_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_5_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_5_A_bx,
      hInputStubs_V_dout     => DL_twoS_5_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_5_A_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_5_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIA_2S_5_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIA_2S_5_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIA_2S_5_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIB_2S_5_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIB_2S_5_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIB_2S_5_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHIC_2S_5_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHIC_2S_5_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHIC_2S_5_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIA_2S_5_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIA_2S_5_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIA_2S_5_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIB_2S_5_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIB_2S_5_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIB_2S_5_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D4PHIC_2S_5_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D4PHIC_2S_5_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D4PHIC_2S_5_A_din,
      hLinkWord_V => "01010000000010000010",
      hPhBnWord_V => "00000000000000000000011100000111"
  );

  LATCH_IR_2S_5_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_5_B_bx,
      start => IR_2S_5_B_start
  );

  IR_2S_5_B : entity work.IR_2S_5_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_5_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_5_B_bx,
      hInputStubs_V_dout     => DL_twoS_5_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_5_B_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_5_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIB_2S_5_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIB_2S_5_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIB_2S_5_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIC_2S_5_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIC_2S_5_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIC_2S_5_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHID_2S_5_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHID_2S_5_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHID_2S_5_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIB_2S_5_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIB_2S_5_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIB_2S_5_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIC_2S_5_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIC_2S_5_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIC_2S_5_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D4PHID_2S_5_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D4PHID_2S_5_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D4PHID_2S_5_B_din,
      hLinkWord_V => "01010000000010000010",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_2S_6_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_6_A_bx,
      start => IR_2S_6_A_start
  );

  IR_2S_6_A : entity work.IR_2S_6_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_6_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_6_A_bx,
      hInputStubs_V_dout     => DL_twoS_6_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_6_A_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_6_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D2PHIA_2S_6_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D2PHIA_2S_6_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D2PHIA_2S_6_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D2PHIB_2S_6_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D2PHIB_2S_6_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D2PHIB_2S_6_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D2PHIC_2S_6_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D2PHIC_2S_6_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D2PHIC_2S_6_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D5PHIA_2S_6_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D5PHIA_2S_6_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D5PHIA_2S_6_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D5PHIB_2S_6_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D5PHIB_2S_6_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D5PHIB_2S_6_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D5PHIC_2S_6_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D5PHIC_2S_6_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D5PHIC_2S_6_A_din,
      hLinkWord_V => "01010000000010100100",
      hPhBnWord_V => "00000000000000000000011100000111"
  );

  LATCH_IR_2S_6_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_2S_6_B_bx,
      start => IR_2S_6_B_start
  );

  IR_2S_6_B : entity work.IR_2S_6_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_2S_6_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_2S_6_B_bx,
      hInputStubs_V_dout     => DL_twoS_6_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_twoS_6_B_link_empty_neg,
      hInputStubs_V_read     => DL_twoS_6_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D2PHIB_2S_6_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D2PHIB_2S_6_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D2PHIB_2S_6_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D2PHIC_2S_6_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D2PHIC_2S_6_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D2PHIC_2S_6_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D2PHID_2S_6_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D2PHID_2S_6_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D2PHID_2S_6_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D5PHIB_2S_6_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D5PHIB_2S_6_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D5PHIB_2S_6_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D5PHIC_2S_6_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D5PHIC_2S_6_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D5PHIC_2S_6_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D5PHID_2S_6_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D5PHID_2S_6_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D5PHID_2S_6_B_din,
      hLinkWord_V => "01010000000010100100",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_neg2S_1_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_1_A_bx,
      start => IR_neg2S_1_A_start
  );

  IR_neg2S_1_A : entity work.IR_neg2S_1_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_1_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_1_A_bx,
      hInputStubs_V_dout     => DL_neg2S_1_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_1_A_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_1_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L4PHIA_neg2S_1_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L4PHIA_neg2S_1_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L4PHIA_neg2S_1_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L4PHIB_neg2S_1_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L4PHIB_neg2S_1_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L4PHIB_neg2S_1_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L4PHIC_neg2S_1_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L4PHIC_neg2S_1_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L4PHIC_neg2S_1_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L5PHIA_neg2S_1_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L5PHIA_neg2S_1_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L5PHIA_neg2S_1_A_din,
      hLinkWord_V => "01010000000010111001",
      hPhBnWord_V => "00000000000000000000000100000111"
  );

  LATCH_IR_neg2S_1_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_1_B_bx,
      start => IR_neg2S_1_B_start
  );

  IR_neg2S_1_B : entity work.IR_neg2S_1_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_1_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_1_B_bx,
      hInputStubs_V_dout     => DL_neg2S_1_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_1_B_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_1_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L4PHIB_neg2S_1_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L4PHIB_neg2S_1_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L4PHIB_neg2S_1_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L4PHIC_neg2S_1_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L4PHIC_neg2S_1_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L4PHIC_neg2S_1_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L4PHID_neg2S_1_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L4PHID_neg2S_1_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L4PHID_neg2S_1_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_L5PHID_neg2S_1_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_L5PHID_neg2S_1_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_L5PHID_neg2S_1_B_din,
      hLinkWord_V => "01010000000010111001",
      hPhBnWord_V => "00000000000000000000100000001110"
  );

  LATCH_IR_neg2S_2_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_2_A_bx,
      start => IR_neg2S_2_A_start
  );

  IR_neg2S_2_A : entity work.IR_neg2S_2_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_2_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_2_A_bx,
      hInputStubs_V_dout     => DL_neg2S_2_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_2_A_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_2_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L5PHIA_neg2S_2_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L5PHIA_neg2S_2_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L5PHIA_neg2S_2_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L5PHIB_neg2S_2_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L5PHIB_neg2S_2_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L5PHIB_neg2S_2_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L5PHIC_neg2S_2_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L5PHIC_neg2S_2_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L5PHIC_neg2S_2_A_din,
      hLinkWord_V => "00110000000000001011",
      hPhBnWord_V => "00000000000000000000000000000111"
  );

  LATCH_IR_neg2S_2_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_2_B_bx,
      start => IR_neg2S_2_B_start
  );

  IR_neg2S_2_B : entity work.IR_neg2S_2_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_2_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_2_B_bx,
      hInputStubs_V_dout     => DL_neg2S_2_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_2_B_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_2_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L5PHIB_neg2S_2_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L5PHIB_neg2S_2_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L5PHIB_neg2S_2_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L5PHIC_neg2S_2_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L5PHIC_neg2S_2_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L5PHIC_neg2S_2_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L5PHID_neg2S_2_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L5PHID_neg2S_2_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L5PHID_neg2S_2_B_din,
      hLinkWord_V => "00110000000000001011",
      hPhBnWord_V => "00000000000000000000000000001110"
  );

  LATCH_IR_neg2S_3_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_3_A_bx,
      start => IR_neg2S_3_A_start
  );

  IR_neg2S_3_A : entity work.IR_neg2S_3_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_3_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_3_A_bx,
      hInputStubs_V_dout     => DL_neg2S_3_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_3_A_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_3_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIA_neg2S_3_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIA_neg2S_3_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIA_neg2S_3_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHIB_neg2S_3_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHIB_neg2S_3_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHIB_neg2S_3_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L6PHIC_neg2S_3_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L6PHIC_neg2S_3_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L6PHIC_neg2S_3_A_din,
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "00000000000000000000000000000111"
  );

  LATCH_IR_neg2S_3_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_3_B_bx,
      start => IR_neg2S_3_B_start
  );

  IR_neg2S_3_B : entity work.IR_neg2S_3_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_3_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_3_B_bx,
      hInputStubs_V_dout     => DL_neg2S_3_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_3_B_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_3_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIC_neg2S_3_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIC_neg2S_3_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIC_neg2S_3_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHID_neg2S_3_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHID_neg2S_3_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHID_neg2S_3_B_din,
      hLinkWord_V => "00110000000000001101",
      hPhBnWord_V => "00000000000000000000000000001100"
  );

  LATCH_IR_neg2S_4_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_4_A_bx,
      start => IR_neg2S_4_A_start
  );

  IR_neg2S_4_A : entity work.IR_neg2S_4_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_4_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_4_A_bx,
      hInputStubs_V_dout     => DL_neg2S_4_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_4_A_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_4_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIA_neg2S_4_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIA_neg2S_4_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIA_neg2S_4_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHIB_neg2S_4_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHIB_neg2S_4_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHIB_neg2S_4_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D3PHIA_neg2S_4_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D3PHIA_neg2S_4_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D3PHIA_neg2S_4_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIB_neg2S_4_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIB_neg2S_4_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIB_neg2S_4_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIC_neg2S_4_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIC_neg2S_4_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIC_neg2S_4_A_din,
      hLinkWord_V => "01010000000001101101",
      hPhBnWord_V => "00000000000000000000011100000011"
  );

  LATCH_IR_neg2S_4_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_4_B_bx,
      start => IR_neg2S_4_B_start
  );

  IR_neg2S_4_B : entity work.IR_neg2S_4_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_4_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_4_B_bx,
      hInputStubs_V_dout     => DL_neg2S_4_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_4_B_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_4_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_L6PHIB_neg2S_4_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_L6PHIB_neg2S_4_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_L6PHIB_neg2S_4_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_L6PHIC_neg2S_4_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_L6PHIC_neg2S_4_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_L6PHIC_neg2S_4_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_L6PHID_neg2S_4_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_L6PHID_neg2S_4_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_L6PHID_neg2S_4_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D3PHIB_neg2S_4_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D3PHIB_neg2S_4_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D3PHIB_neg2S_4_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D3PHIC_neg2S_4_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D3PHIC_neg2S_4_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D3PHIC_neg2S_4_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D3PHID_neg2S_4_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D3PHID_neg2S_4_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D3PHID_neg2S_4_B_din,
      hLinkWord_V => "01010000000001101101",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_neg2S_5_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_5_A_bx,
      start => IR_neg2S_5_A_start
  );

  IR_neg2S_5_A : entity work.IR_neg2S_5_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_5_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_5_A_bx,
      hInputStubs_V_dout     => DL_neg2S_5_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_5_A_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_5_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIA_neg2S_5_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIA_neg2S_5_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIA_neg2S_5_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIB_neg2S_5_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIB_neg2S_5_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIB_neg2S_5_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHIC_neg2S_5_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHIC_neg2S_5_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHIC_neg2S_5_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIA_neg2S_5_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIA_neg2S_5_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIA_neg2S_5_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIB_neg2S_5_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIB_neg2S_5_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIB_neg2S_5_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D4PHIC_neg2S_5_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D4PHIC_neg2S_5_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D4PHIC_neg2S_5_A_din,
      hLinkWord_V => "01010000000010000010",
      hPhBnWord_V => "00000000000000000000011100000111"
  );

  LATCH_IR_neg2S_5_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_5_B_bx,
      start => IR_neg2S_5_B_start
  );

  IR_neg2S_5_B : entity work.IR_neg2S_5_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_5_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_5_B_bx,
      hInputStubs_V_dout     => DL_neg2S_5_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_5_B_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_5_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D1PHIB_neg2S_5_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D1PHIB_neg2S_5_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D1PHIB_neg2S_5_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D1PHIC_neg2S_5_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D1PHIC_neg2S_5_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D1PHIC_neg2S_5_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D1PHID_neg2S_5_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D1PHID_neg2S_5_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D1PHID_neg2S_5_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D4PHIB_neg2S_5_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D4PHIB_neg2S_5_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D4PHIB_neg2S_5_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D4PHIC_neg2S_5_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D4PHIC_neg2S_5_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D4PHIC_neg2S_5_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D4PHID_neg2S_5_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D4PHID_neg2S_5_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D4PHID_neg2S_5_B_din,
      hLinkWord_V => "01010000000010000010",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_IR_neg2S_6_A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_6_A_bx,
      start => IR_neg2S_6_A_start
  );

  IR_neg2S_6_A : entity work.IR_neg2S_6_A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_6_A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_6_A_bx,
      hInputStubs_V_dout     => DL_neg2S_6_A_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_6_A_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_6_A_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D2PHIA_neg2S_6_A_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D2PHIA_neg2S_6_A_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D2PHIA_neg2S_6_A_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D2PHIB_neg2S_6_A_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D2PHIB_neg2S_6_A_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D2PHIB_neg2S_6_A_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D2PHIC_neg2S_6_A_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D2PHIC_neg2S_6_A_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D2PHIC_neg2S_6_A_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D5PHIA_neg2S_6_A_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D5PHIA_neg2S_6_A_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D5PHIA_neg2S_6_A_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D5PHIB_neg2S_6_A_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D5PHIB_neg2S_6_A_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D5PHIB_neg2S_6_A_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D5PHIC_neg2S_6_A_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D5PHIC_neg2S_6_A_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D5PHIC_neg2S_6_A_din,
      hLinkWord_V => "01010000000010100100",
      hPhBnWord_V => "00000000000000000000011100000111"
  );

  LATCH_IR_neg2S_6_B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_start,
      bx_out => IR_bx_in,
      bx => IR_neg2S_6_B_bx,
      start => IR_neg2S_6_B_start
  );

  IR_neg2S_6_B : entity work.IR_neg2S_6_B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => IR_neg2S_6_B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => IR_neg2S_6_B_bx,
      hInputStubs_V_dout     => DL_neg2S_6_B_link_AV_dout,
      hInputStubs_V_empty_n  => DL_neg2S_6_B_link_empty_neg,
      hInputStubs_V_read     => DL_neg2S_6_B_link_read,
      hOutputStubs_0_dataarray_data_V_ce0       => open,
      hOutputStubs_0_dataarray_data_V_we0       => IL_D2PHIB_neg2S_6_B_wea,
      hOutputStubs_0_dataarray_data_V_address0  => IL_D2PHIB_neg2S_6_B_writeaddr,
      hOutputStubs_0_dataarray_data_V_d0        => IL_D2PHIB_neg2S_6_B_din,
      hOutputStubs_1_dataarray_data_V_ce0       => open,
      hOutputStubs_1_dataarray_data_V_we0       => IL_D2PHIC_neg2S_6_B_wea,
      hOutputStubs_1_dataarray_data_V_address0  => IL_D2PHIC_neg2S_6_B_writeaddr,
      hOutputStubs_1_dataarray_data_V_d0        => IL_D2PHIC_neg2S_6_B_din,
      hOutputStubs_2_dataarray_data_V_ce0       => open,
      hOutputStubs_2_dataarray_data_V_we0       => IL_D2PHID_neg2S_6_B_wea,
      hOutputStubs_2_dataarray_data_V_address0  => IL_D2PHID_neg2S_6_B_writeaddr,
      hOutputStubs_2_dataarray_data_V_d0        => IL_D2PHID_neg2S_6_B_din,
      hOutputStubs_3_dataarray_data_V_ce0       => open,
      hOutputStubs_3_dataarray_data_V_we0       => IL_D5PHIB_neg2S_6_B_wea,
      hOutputStubs_3_dataarray_data_V_address0  => IL_D5PHIB_neg2S_6_B_writeaddr,
      hOutputStubs_3_dataarray_data_V_d0        => IL_D5PHIB_neg2S_6_B_din,
      hOutputStubs_4_dataarray_data_V_ce0       => open,
      hOutputStubs_4_dataarray_data_V_we0       => IL_D5PHIC_neg2S_6_B_wea,
      hOutputStubs_4_dataarray_data_V_address0  => IL_D5PHIC_neg2S_6_B_writeaddr,
      hOutputStubs_4_dataarray_data_V_d0        => IL_D5PHIC_neg2S_6_B_din,
      hOutputStubs_5_dataarray_data_V_ce0       => open,
      hOutputStubs_5_dataarray_data_V_we0       => IL_D5PHID_neg2S_6_B_wea,
      hOutputStubs_5_dataarray_data_V_address0  => IL_D5PHID_neg2S_6_B_writeaddr,
      hOutputStubs_5_dataarray_data_V_d0        => IL_D5PHID_neg2S_6_B_din,
      hLinkWord_V => "01010000000010100100",
      hPhBnWord_V => "00000000000000000000111000001110"
  );

  LATCH_VMR_L1PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHIA_bx,
      start => VMR_L1PHIA_start
  );

  VMR_L1PHIA : entity work.VMR_L1PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => VMR_done,
      bx_V          => VMR_L1PHIA_bx,
      bx_o_V        => VMR_bx_out,
      bx_o_V_ap_vld => open,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHIA_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHIA_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHIA_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHIA_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHIA_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHIA_PS10G_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHIA_PS10G_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHIA_PS10G_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHIA_PS10G_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHIA_PS10G_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHIA_negPS10G_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHIA_negPS10G_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHIA_negPS10G_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHIA_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHIA_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L1PHIA_negPS10G_2_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L1PHIA_negPS10G_2_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L1PHIA_negPS10G_2_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L1PHIA_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L1PHIA_negPS10G_2_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIAn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHIA_BF_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHIA_BF_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHIA_BF_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHIA_BE_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHIA_BE_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHIA_BE_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHIA_OM_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHIA_OM_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHIA_OM_din
  );

  LATCH_VMR_L1PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHIB_bx,
      start => VMR_L1PHIB_start
  );

  VMR_L1PHIB : entity work.VMR_L1PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L1PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHIB_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHIB_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHIB_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHIB_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHIB_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHIB_PS10G_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHIB_PS10G_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHIB_PS10G_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHIB_PS10G_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHIB_PS10G_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHIB_negPS10G_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHIB_negPS10G_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHIB_negPS10G_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHIB_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHIB_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L1PHIB_negPS10G_2_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L1PHIB_negPS10G_2_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L1PHIB_negPS10G_2_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L1PHIB_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L1PHIB_negPS10G_2_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIBn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHIB_BD_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHIB_BD_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHIB_BD_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHIB_BC_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHIB_BC_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHIB_BC_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHIB_BA_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHIB_BA_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHIB_BA_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L1PHIB_OM_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L1PHIB_OM_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L1PHIB_OM_din,
      memoriesASInner_4_dataarray_data_V_ce0       => open,
      memoriesASInner_4_dataarray_data_V_we0       => AS_L1PHIB_OR_wea,
      memoriesASInner_4_dataarray_data_V_address0  => AS_L1PHIB_OR_writeaddr,
      memoriesASInner_4_dataarray_data_V_d0        => AS_L1PHIB_OR_din
  );

  LATCH_VMR_L1PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHIC_bx,
      start => VMR_L1PHIC_start
  );

  VMR_L1PHIC : entity work.VMR_L1PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L1PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHIC_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHIC_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHIC_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHIC_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHIC_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHIC_PS10G_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHIC_PS10G_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHIC_PS10G_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHIC_PS10G_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHIC_PS10G_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHIC_negPS10G_2_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHIC_negPS10G_2_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHIC_negPS10G_2_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHIC_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHIC_negPS10G_2_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHICn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHIC_BB_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHIC_BB_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHIC_BB_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHIC_BF_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHIC_BF_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHIC_BF_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHIC_BE_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHIC_BE_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHIC_BE_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L1PHIC_OL_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L1PHIC_OL_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L1PHIC_OL_din,
      memoriesASInner_4_dataarray_data_V_ce0       => open,
      memoriesASInner_4_dataarray_data_V_we0       => AS_L1PHIC_OM_wea,
      memoriesASInner_4_dataarray_data_V_address0  => AS_L1PHIC_OM_writeaddr,
      memoriesASInner_4_dataarray_data_V_d0        => AS_L1PHIC_OM_din
  );

  LATCH_VMR_L1PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHID_bx,
      start => VMR_L1PHID_start
  );

  VMR_L1PHID : entity work.VMR_L1PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L1PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHID_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHID_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHID_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHID_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHID_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHID_PS10G_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHID_PS10G_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHID_PS10G_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHID_PS10G_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHID_PS10G_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHID_PS10G_2_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHID_PS10G_2_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHID_PS10G_2_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHID_PS10G_2_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHID_PS10G_2_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L1PHID_negPS10G_1_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L1PHID_negPS10G_1_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L1PHID_negPS10G_1_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L1PHID_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L1PHID_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_L1PHID_negPS10G_2_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_L1PHID_negPS10G_2_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_L1PHID_negPS10G_2_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_L1PHID_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_L1PHID_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_L1PHID_negPS10G_2_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_L1PHID_negPS10G_2_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_L1PHID_negPS10G_2_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_L1PHID_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_L1PHID_negPS10G_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIDn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHID_BD_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHID_BD_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHID_BD_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHID_BC_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHID_BC_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHID_BC_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHID_BA_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHID_BA_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHID_BA_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L1PHID_OM_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L1PHID_OM_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L1PHID_OM_din,
      memoriesASInner_4_dataarray_data_V_ce0       => open,
      memoriesASInner_4_dataarray_data_V_we0       => AS_L1PHID_OR_wea,
      memoriesASInner_4_dataarray_data_V_address0  => AS_L1PHID_OR_writeaddr,
      memoriesASInner_4_dataarray_data_V_d0        => AS_L1PHID_OR_din
  );

  LATCH_VMR_L1PHIE: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHIE_bx,
      start => VMR_L1PHIE_start
  );

  VMR_L1PHIE : entity work.VMR_L1PHIE
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHIE_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L1PHIE_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHIE_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHIE_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHIE_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHIE_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHIE_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHIE_PS10G_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHIE_PS10G_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHIE_PS10G_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHIE_PS10G_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHIE_PS10G_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHIE_PS10G_2_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHIE_PS10G_2_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHIE_PS10G_2_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHIE_PS10G_2_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHIE_PS10G_2_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L1PHIE_negPS10G_1_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L1PHIE_negPS10G_1_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L1PHIE_negPS10G_1_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L1PHIE_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L1PHIE_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_L1PHIE_negPS10G_2_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_L1PHIE_negPS10G_2_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_L1PHIE_negPS10G_2_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_L1PHIE_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_L1PHIE_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_L1PHIE_negPS10G_2_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_L1PHIE_negPS10G_2_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_L1PHIE_negPS10G_2_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_L1PHIE_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_L1PHIE_negPS10G_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIEn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIEn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIEn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHIE_BB_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHIE_BB_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHIE_BB_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHIE_BF_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHIE_BF_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHIE_BF_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHIE_BE_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHIE_BE_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHIE_BE_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L1PHIE_OL_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L1PHIE_OL_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L1PHIE_OL_din,
      memoriesASInner_4_dataarray_data_V_ce0       => open,
      memoriesASInner_4_dataarray_data_V_we0       => AS_L1PHIE_OM_wea,
      memoriesASInner_4_dataarray_data_V_address0  => AS_L1PHIE_OM_writeaddr,
      memoriesASInner_4_dataarray_data_V_d0        => AS_L1PHIE_OM_din
  );

  LATCH_VMR_L1PHIF: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHIF_bx,
      start => VMR_L1PHIF_start
  );

  VMR_L1PHIF : entity work.VMR_L1PHIF
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHIF_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L1PHIF_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHIF_PS10G_2_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHIF_PS10G_2_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHIF_PS10G_2_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHIF_PS10G_2_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHIF_PS10G_2_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHIF_negPS10G_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHIF_negPS10G_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHIF_negPS10G_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHIF_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHIF_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHIF_negPS10G_2_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHIF_negPS10G_2_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHIF_negPS10G_2_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHIF_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHIF_negPS10G_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIFn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIFn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIFn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHIF_BD_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHIF_BD_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHIF_BD_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHIF_BC_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHIF_BC_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHIF_BC_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHIF_BA_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHIF_BA_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHIF_BA_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L1PHIF_OM_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L1PHIF_OM_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L1PHIF_OM_din,
      memoriesASInner_4_dataarray_data_V_ce0       => open,
      memoriesASInner_4_dataarray_data_V_we0       => AS_L1PHIF_OR_wea,
      memoriesASInner_4_dataarray_data_V_address0  => AS_L1PHIF_OR_writeaddr,
      memoriesASInner_4_dataarray_data_V_d0        => AS_L1PHIF_OR_din
  );

  LATCH_VMR_L1PHIG: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHIG_bx,
      start => VMR_L1PHIG_start
  );

  VMR_L1PHIG : entity work.VMR_L1PHIG
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHIG_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L1PHIG_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHIG_PS10G_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHIG_PS10G_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHIG_PS10G_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHIG_PS10G_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHIG_PS10G_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHIG_PS10G_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHIG_PS10G_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHIG_PS10G_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHIG_PS10G_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHIG_PS10G_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHIG_negPS10G_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHIG_negPS10G_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHIG_negPS10G_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHIG_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHIG_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L1PHIG_negPS10G_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L1PHIG_negPS10G_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L1PHIG_negPS10G_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L1PHIG_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L1PHIG_negPS10G_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIGn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIGn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIGn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHIG_BB_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHIG_BB_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHIG_BB_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHIG_BF_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHIG_BF_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHIG_BF_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHIG_BE_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHIG_BE_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHIG_BE_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L1PHIG_OL_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L1PHIG_OL_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L1PHIG_OL_din,
      memoriesASInner_4_dataarray_data_V_ce0       => open,
      memoriesASInner_4_dataarray_data_V_we0       => AS_L1PHIG_OM_wea,
      memoriesASInner_4_dataarray_data_V_address0  => AS_L1PHIG_OM_writeaddr,
      memoriesASInner_4_dataarray_data_V_d0        => AS_L1PHIG_OM_din
  );

  LATCH_VMR_L1PHIH: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L1PHIH_bx,
      start => VMR_L1PHIH_start
  );

  VMR_L1PHIH : entity work.VMR_L1PHIH
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L1PHIH_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L1PHIH_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L1PHIH_PS10G_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L1PHIH_PS10G_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L1PHIH_PS10G_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L1PHIH_PS10G_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L1PHIH_PS10G_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L1PHIH_PS10G_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L1PHIH_PS10G_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L1PHIH_PS10G_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L1PHIH_PS10G_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L1PHIH_PS10G_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L1PHIH_negPS10G_2_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L1PHIH_negPS10G_2_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L1PHIH_negPS10G_2_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L1PHIH_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L1PHIH_negPS10G_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L1PHIHn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L1PHIHn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L1PHIHn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L1PHIH_BD_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L1PHIH_BD_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L1PHIH_BD_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L1PHIH_BC_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L1PHIH_BC_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L1PHIH_BC_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L1PHIH_OM_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L1PHIH_OM_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L1PHIH_OM_din
  );

  LATCH_VMR_L2PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L2PHIA_bx,
      start => VMR_L2PHIA_start
  );

  VMR_L2PHIA : entity work.VMR_L2PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L2PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L2PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L2PHIA_PS10G_3_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L2PHIA_PS10G_3_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L2PHIA_PS10G_3_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L2PHIA_PS10G_3_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L2PHIA_PS10G_3_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L2PHIA_negPS10G_3_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L2PHIA_negPS10G_3_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L2PHIA_negPS10G_3_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L2PHIA_negPS10G_3_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L2PHIA_negPS10G_3_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHIAn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L2PHIA_B_L1A_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L2PHIA_B_L1A_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L2PHIA_B_L1A_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_L2PHIA_B_L1B_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_L2PHIA_B_L1B_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_L2PHIA_B_L1B_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_L2PHIA_B_L1C_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_L2PHIA_B_L1C_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_L2PHIA_B_L1C_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L2PHIA_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L2PHIA_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L2PHIA_BM_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L2PHIA_OM_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L2PHIA_OM_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L2PHIA_OM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L2PHIAn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L2PHIAn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L2PHIAn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_L2PHIAn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_L2PHIAn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_L2PHIAn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_L2PHIAn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_L2PHIAn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_L2PHIAn3_din
  );

  LATCH_VMR_L2PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L2PHIB_bx,
      start => VMR_L2PHIB_start
  );

  VMR_L2PHIB : entity work.VMR_L2PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L2PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L2PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L2PHIB_PS10G_3_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L2PHIB_PS10G_3_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L2PHIB_PS10G_3_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L2PHIB_PS10G_3_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L2PHIB_PS10G_3_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L2PHIB_PS10G_3_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L2PHIB_PS10G_3_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L2PHIB_PS10G_3_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L2PHIB_PS10G_3_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L2PHIB_PS10G_3_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L2PHIB_negPS10G_3_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L2PHIB_negPS10G_3_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L2PHIB_negPS10G_3_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L2PHIB_negPS10G_3_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L2PHIB_negPS10G_3_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L2PHIB_negPS10G_3_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L2PHIB_negPS10G_3_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L2PHIB_negPS10G_3_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L2PHIB_negPS10G_3_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L2PHIB_negPS10G_3_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHIBn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L2PHIB_B_L1D_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L2PHIB_B_L1D_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L2PHIB_B_L1D_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_L2PHIB_B_L1E_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_L2PHIB_B_L1E_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_L2PHIB_B_L1E_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_L2PHIB_B_L1F_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_L2PHIB_B_L1F_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_L2PHIB_B_L1F_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L2PHIB_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L2PHIB_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L2PHIB_BM_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L2PHIB_BR_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L2PHIB_BR_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L2PHIB_BR_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L2PHIB_OM_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L2PHIB_OM_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L2PHIB_OM_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L2PHIB_OR_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L2PHIB_OR_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L2PHIB_OR_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L2PHIBn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L2PHIBn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L2PHIBn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_L2PHIBn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_L2PHIBn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_L2PHIBn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_L2PHIBn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_L2PHIBn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_L2PHIBn3_din
  );

  LATCH_VMR_L2PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L2PHIC_bx,
      start => VMR_L2PHIC_start
  );

  VMR_L2PHIC : entity work.VMR_L2PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L2PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L2PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L2PHIC_PS10G_3_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L2PHIC_PS10G_3_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L2PHIC_PS10G_3_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L2PHIC_PS10G_3_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L2PHIC_PS10G_3_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L2PHIC_PS10G_3_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L2PHIC_PS10G_3_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L2PHIC_PS10G_3_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L2PHIC_PS10G_3_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L2PHIC_PS10G_3_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L2PHIC_negPS10G_3_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L2PHIC_negPS10G_3_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L2PHIC_negPS10G_3_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L2PHIC_negPS10G_3_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L2PHIC_negPS10G_3_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L2PHIC_negPS10G_3_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L2PHIC_negPS10G_3_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L2PHIC_negPS10G_3_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L2PHIC_negPS10G_3_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L2PHIC_negPS10G_3_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHICn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L2PHIC_B_L1G_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L2PHIC_B_L1G_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L2PHIC_B_L1G_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_L2PHIC_B_L1H_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_L2PHIC_B_L1H_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_L2PHIC_B_L1H_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_L2PHIC_B_L1I_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_L2PHIC_B_L1I_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_L2PHIC_B_L1I_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L2PHIC_BL_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L2PHIC_BL_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L2PHIC_BL_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L2PHIC_BM_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L2PHIC_BM_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L2PHIC_BM_din,
      memoriesASInner_2_dataarray_data_V_ce0       => open,
      memoriesASInner_2_dataarray_data_V_we0       => AS_L2PHIC_OL_wea,
      memoriesASInner_2_dataarray_data_V_address0  => AS_L2PHIC_OL_writeaddr,
      memoriesASInner_2_dataarray_data_V_d0        => AS_L2PHIC_OL_din,
      memoriesASInner_3_dataarray_data_V_ce0       => open,
      memoriesASInner_3_dataarray_data_V_we0       => AS_L2PHIC_OM_wea,
      memoriesASInner_3_dataarray_data_V_address0  => AS_L2PHIC_OM_writeaddr,
      memoriesASInner_3_dataarray_data_V_d0        => AS_L2PHIC_OM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L2PHICn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L2PHICn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L2PHICn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_L2PHICn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_L2PHICn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_L2PHICn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_L2PHICn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_L2PHICn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_L2PHICn3_din
  );

  LATCH_VMR_L2PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L2PHID_bx,
      start => VMR_L2PHID_start
  );

  VMR_L2PHID : entity work.VMR_L2PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L2PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L2PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L2PHID_PS10G_3_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L2PHID_PS10G_3_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L2PHID_PS10G_3_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L2PHID_PS10G_3_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L2PHID_PS10G_3_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L2PHID_negPS10G_3_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L2PHID_negPS10G_3_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L2PHID_negPS10G_3_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L2PHID_negPS10G_3_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L2PHID_negPS10G_3_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L2PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L2PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L2PHIDn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L2PHID_B_L1J_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L2PHID_B_L1J_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L2PHID_B_L1J_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_L2PHID_B_L1K_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_L2PHID_B_L1K_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_L2PHID_B_L1K_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_L2PHID_B_L1L_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_L2PHID_B_L1L_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_L2PHID_B_L1L_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L2PHID_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L2PHID_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L2PHID_BM_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L2PHID_OM_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L2PHID_OM_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L2PHID_OM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L2PHIDn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L2PHIDn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L2PHIDn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_L2PHIDn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_L2PHIDn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_L2PHIDn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_L2PHIDn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_L2PHIDn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_L2PHIDn3_din
  );

  LATCH_VMR_L3PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L3PHIA_bx,
      start => VMR_L3PHIA_start
  );

  VMR_L3PHIA : entity work.VMR_L3PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L3PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L3PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L3PHIA_PS_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L3PHIA_PS_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L3PHIA_PS_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L3PHIA_PS_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L3PHIA_PS_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L3PHIA_PS_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L3PHIA_PS_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L3PHIA_PS_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L3PHIA_PS_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L3PHIA_PS_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L3PHIA_negPS_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L3PHIA_negPS_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L3PHIA_negPS_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L3PHIA_negPS_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L3PHIA_negPS_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L3PHIA_negPS_2_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L3PHIA_negPS_2_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L3PHIA_negPS_2_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L3PHIA_negPS_2_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L3PHIA_negPS_2_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHIAn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L3PHIA_B_L2A_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L3PHIA_B_L2A_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L3PHIA_B_L2A_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L3PHIA_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L3PHIA_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L3PHIA_BM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L3PHIIn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L3PHIIn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L3PHIIn1_din
  );

  LATCH_VMR_L3PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L3PHIB_bx,
      start => VMR_L3PHIB_start
  );

  VMR_L3PHIB : entity work.VMR_L3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L3PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L3PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L3PHIB_PS_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L3PHIB_PS_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L3PHIB_PS_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L3PHIB_PS_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L3PHIB_PS_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L3PHIB_PS_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L3PHIB_PS_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L3PHIB_PS_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L3PHIB_PS_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L3PHIB_PS_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L3PHIB_PS_2_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L3PHIB_PS_2_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L3PHIB_PS_2_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L3PHIB_PS_2_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L3PHIB_PS_2_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L3PHIB_negPS_1_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L3PHIB_negPS_1_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L3PHIB_negPS_1_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L3PHIB_negPS_1_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L3PHIB_negPS_1_A_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_L3PHIB_negPS_1_B_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_L3PHIB_negPS_1_B_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_L3PHIB_negPS_1_B_V_dout,
      inputStubs_4_nentries_0_V               => IL_L3PHIB_negPS_1_B_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_L3PHIB_negPS_1_B_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_L3PHIB_negPS_2_A_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_L3PHIB_negPS_2_A_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_L3PHIB_negPS_2_A_V_dout,
      inputStubs_5_nentries_0_V               => IL_L3PHIB_negPS_2_A_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_L3PHIB_negPS_2_A_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_L3PHIB_negPS_2_B_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_L3PHIB_negPS_2_B_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_L3PHIB_negPS_2_B_V_dout,
      inputStubs_6_nentries_0_V               => IL_L3PHIB_negPS_2_B_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_L3PHIB_negPS_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHIBn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L3PHIB_B_L2B_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L3PHIB_B_L2B_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L3PHIB_B_L2B_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L3PHIB_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L3PHIB_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L3PHIB_BM_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L3PHIB_BR_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L3PHIB_BR_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L3PHIB_BR_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L3PHIJn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L3PHIJn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L3PHIJn1_din
  );

  LATCH_VMR_L3PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L3PHIC_bx,
      start => VMR_L3PHIC_start
  );

  VMR_L3PHIC : entity work.VMR_L3PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L3PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L3PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L3PHIC_PS_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L3PHIC_PS_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L3PHIC_PS_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L3PHIC_PS_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L3PHIC_PS_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L3PHIC_PS_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L3PHIC_PS_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L3PHIC_PS_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L3PHIC_PS_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L3PHIC_PS_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L3PHIC_negPS_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L3PHIC_negPS_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L3PHIC_negPS_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L3PHIC_negPS_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L3PHIC_negPS_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L3PHIC_negPS_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L3PHIC_negPS_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L3PHIC_negPS_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L3PHIC_negPS_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L3PHIC_negPS_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHICn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L3PHIC_B_L2C_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L3PHIC_B_L2C_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L3PHIC_B_L2C_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L3PHIC_BL_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L3PHIC_BL_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L3PHIC_BL_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L3PHIC_BM_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L3PHIC_BM_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L3PHIC_BM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L3PHIKn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L3PHIKn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L3PHIKn1_din
  );

  LATCH_VMR_L3PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L3PHID_bx,
      start => VMR_L3PHID_start
  );

  VMR_L3PHID : entity work.VMR_L3PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L3PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L3PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L3PHID_PS_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L3PHID_PS_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L3PHID_PS_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L3PHID_PS_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L3PHID_PS_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L3PHID_PS_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L3PHID_PS_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L3PHID_PS_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L3PHID_PS_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L3PHID_PS_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L3PHID_negPS_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L3PHID_negPS_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L3PHID_negPS_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L3PHID_negPS_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L3PHID_negPS_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L3PHID_negPS_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L3PHID_negPS_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L3PHID_negPS_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L3PHID_negPS_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L3PHID_negPS_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L3PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L3PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L3PHIDn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L3PHID_B_L2D_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L3PHID_B_L2D_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L3PHID_B_L2D_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L3PHID_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L3PHID_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L3PHID_BM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L3PHILn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L3PHILn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L3PHILn1_din
  );

  LATCH_VMR_L4PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L4PHIA_bx,
      start => VMR_L4PHIA_start
  );

  VMR_L4PHIA : entity work.VMR_L4PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L4PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L4PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L4PHIA_2S_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L4PHIA_2S_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L4PHIA_2S_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L4PHIA_2S_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L4PHIA_2S_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L4PHIA_neg2S_1_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L4PHIA_neg2S_1_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L4PHIA_neg2S_1_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L4PHIA_neg2S_1_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L4PHIA_neg2S_1_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHIAn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L4PHIA_B_L3A_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L4PHIA_B_L3A_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L4PHIA_B_L3A_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L4PHIAn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L4PHIAn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L4PHIAn1_din
  );

  LATCH_VMR_L4PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L4PHIB_bx,
      start => VMR_L4PHIB_start
  );

  VMR_L4PHIB : entity work.VMR_L4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L4PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L4PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L4PHIB_2S_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L4PHIB_2S_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L4PHIB_2S_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L4PHIB_2S_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L4PHIB_2S_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L4PHIB_2S_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L4PHIB_2S_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L4PHIB_2S_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L4PHIB_2S_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L4PHIB_2S_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L4PHIB_neg2S_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L4PHIB_neg2S_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L4PHIB_neg2S_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L4PHIB_neg2S_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L4PHIB_neg2S_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L4PHIB_neg2S_1_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L4PHIB_neg2S_1_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L4PHIB_neg2S_1_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L4PHIB_neg2S_1_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L4PHIB_neg2S_1_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHIBn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L4PHIB_B_L3B_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L4PHIB_B_L3B_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L4PHIB_B_L3B_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L4PHIBn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L4PHIBn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L4PHIBn1_din
  );

  LATCH_VMR_L4PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L4PHIC_bx,
      start => VMR_L4PHIC_start
  );

  VMR_L4PHIC : entity work.VMR_L4PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L4PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L4PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L4PHIC_2S_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L4PHIC_2S_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L4PHIC_2S_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L4PHIC_2S_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L4PHIC_2S_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L4PHIC_2S_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L4PHIC_2S_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L4PHIC_2S_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L4PHIC_2S_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L4PHIC_2S_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L4PHIC_neg2S_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L4PHIC_neg2S_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L4PHIC_neg2S_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L4PHIC_neg2S_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L4PHIC_neg2S_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L4PHIC_neg2S_1_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L4PHIC_neg2S_1_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L4PHIC_neg2S_1_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L4PHIC_neg2S_1_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L4PHIC_neg2S_1_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHICn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L4PHIC_B_L3C_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L4PHIC_B_L3C_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L4PHIC_B_L3C_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L4PHICn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L4PHICn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L4PHICn1_din
  );

  LATCH_VMR_L4PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L4PHID_bx,
      start => VMR_L4PHID_start
  );

  VMR_L4PHID : entity work.VMR_L4PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L4PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L4PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L4PHID_2S_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L4PHID_2S_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L4PHID_2S_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L4PHID_2S_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L4PHID_2S_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L4PHID_neg2S_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L4PHID_neg2S_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L4PHID_neg2S_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L4PHID_neg2S_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L4PHID_neg2S_1_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L4PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L4PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L4PHIDn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L4PHID_B_L3D_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L4PHID_B_L3D_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L4PHID_B_L3D_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L4PHIDn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L4PHIDn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L4PHIDn1_din
  );

  LATCH_VMR_L5PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L5PHIA_bx,
      start => VMR_L5PHIA_start
  );

  VMR_L5PHIA : entity work.VMR_L5PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L5PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L5PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L5PHIA_2S_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L5PHIA_2S_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L5PHIA_2S_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L5PHIA_2S_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L5PHIA_2S_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L5PHIA_2S_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L5PHIA_2S_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L5PHIA_2S_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L5PHIA_2S_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L5PHIA_2S_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L5PHIA_neg2S_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L5PHIA_neg2S_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L5PHIA_neg2S_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L5PHIA_neg2S_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L5PHIA_neg2S_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L5PHIA_neg2S_2_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L5PHIA_neg2S_2_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L5PHIA_neg2S_2_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L5PHIA_neg2S_2_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L5PHIA_neg2S_2_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHIAn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L5PHIA_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L5PHIA_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L5PHIA_BM_din
  );

  LATCH_VMR_L5PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L5PHIB_bx,
      start => VMR_L5PHIB_start
  );

  VMR_L5PHIB : entity work.VMR_L5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L5PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L5PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L5PHIB_2S_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L5PHIB_2S_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L5PHIB_2S_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L5PHIB_2S_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L5PHIB_2S_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L5PHIB_2S_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L5PHIB_2S_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L5PHIB_2S_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L5PHIB_2S_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L5PHIB_2S_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L5PHIB_neg2S_2_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L5PHIB_neg2S_2_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L5PHIB_neg2S_2_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L5PHIB_neg2S_2_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L5PHIB_neg2S_2_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L5PHIB_neg2S_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L5PHIB_neg2S_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L5PHIB_neg2S_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L5PHIB_neg2S_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L5PHIB_neg2S_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHIBn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L5PHIB_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L5PHIB_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L5PHIB_BM_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L5PHIB_BR_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L5PHIB_BR_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L5PHIB_BR_din
  );

  LATCH_VMR_L5PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L5PHIC_bx,
      start => VMR_L5PHIC_start
  );

  VMR_L5PHIC : entity work.VMR_L5PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L5PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L5PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L5PHIC_2S_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L5PHIC_2S_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L5PHIC_2S_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L5PHIC_2S_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L5PHIC_2S_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L5PHIC_2S_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L5PHIC_2S_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L5PHIC_2S_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L5PHIC_2S_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L5PHIC_2S_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L5PHIC_neg2S_2_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L5PHIC_neg2S_2_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L5PHIC_neg2S_2_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L5PHIC_neg2S_2_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L5PHIC_neg2S_2_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L5PHIC_neg2S_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L5PHIC_neg2S_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L5PHIC_neg2S_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L5PHIC_neg2S_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L5PHIC_neg2S_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHICn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L5PHIC_BL_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L5PHIC_BL_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L5PHIC_BL_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_L5PHIC_BM_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_L5PHIC_BM_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_L5PHIC_BM_din
  );

  LATCH_VMR_L5PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L5PHID_bx,
      start => VMR_L5PHID_start
  );

  VMR_L5PHID : entity work.VMR_L5PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L5PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L5PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L5PHID_2S_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L5PHID_2S_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L5PHID_2S_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L5PHID_2S_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L5PHID_2S_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L5PHID_2S_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L5PHID_2S_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L5PHID_2S_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L5PHID_2S_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L5PHID_2S_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L5PHID_neg2S_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L5PHID_neg2S_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L5PHID_neg2S_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L5PHID_neg2S_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L5PHID_neg2S_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L5PHID_neg2S_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L5PHID_neg2S_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L5PHID_neg2S_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L5PHID_neg2S_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L5PHID_neg2S_2_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L5PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L5PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L5PHIDn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_L5PHID_BM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_L5PHID_BM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_L5PHID_BM_din
  );

  LATCH_VMR_L6PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L6PHIA_bx,
      start => VMR_L6PHIA_start
  );

  VMR_L6PHIA : entity work.VMR_L6PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L6PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L6PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L6PHIA_2S_3_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L6PHIA_2S_3_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L6PHIA_2S_3_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L6PHIA_2S_3_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L6PHIA_2S_3_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L6PHIA_2S_4_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L6PHIA_2S_4_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L6PHIA_2S_4_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L6PHIA_2S_4_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L6PHIA_2S_4_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L6PHIA_neg2S_3_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L6PHIA_neg2S_3_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L6PHIA_neg2S_3_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_L6PHIA_neg2S_3_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L6PHIA_neg2S_3_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L6PHIA_neg2S_4_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L6PHIA_neg2S_4_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L6PHIA_neg2S_4_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L6PHIA_neg2S_4_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L6PHIA_neg2S_4_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHIAn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L6PHIA_B_L5A_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L6PHIA_B_L5A_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L6PHIA_B_L5A_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L6PHIAn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L6PHIAn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L6PHIAn1_din
  );

  LATCH_VMR_L6PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L6PHIB_bx,
      start => VMR_L6PHIB_start
  );

  VMR_L6PHIB : entity work.VMR_L6PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L6PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L6PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L6PHIB_2S_3_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L6PHIB_2S_3_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L6PHIB_2S_3_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L6PHIB_2S_3_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L6PHIB_2S_3_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L6PHIB_2S_4_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L6PHIB_2S_4_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L6PHIB_2S_4_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_L6PHIB_2S_4_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L6PHIB_2S_4_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L6PHIB_2S_4_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L6PHIB_2S_4_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L6PHIB_2S_4_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L6PHIB_2S_4_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L6PHIB_2S_4_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L6PHIB_neg2S_3_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L6PHIB_neg2S_3_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L6PHIB_neg2S_3_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L6PHIB_neg2S_3_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L6PHIB_neg2S_3_A_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_L6PHIB_neg2S_4_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_L6PHIB_neg2S_4_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_L6PHIB_neg2S_4_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_L6PHIB_neg2S_4_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_L6PHIB_neg2S_4_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_L6PHIB_neg2S_4_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_L6PHIB_neg2S_4_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_L6PHIB_neg2S_4_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_L6PHIB_neg2S_4_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_L6PHIB_neg2S_4_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHIBn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L6PHIB_B_L5B_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L6PHIB_B_L5B_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L6PHIB_B_L5B_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L6PHIBn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L6PHIBn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L6PHIBn1_din
  );

  LATCH_VMR_L6PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L6PHIC_bx,
      start => VMR_L6PHIC_start
  );

  VMR_L6PHIC : entity work.VMR_L6PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L6PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L6PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L6PHIC_2S_3_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L6PHIC_2S_3_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L6PHIC_2S_3_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_L6PHIC_2S_3_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L6PHIC_2S_3_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L6PHIC_2S_3_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L6PHIC_2S_3_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L6PHIC_2S_3_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L6PHIC_2S_3_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L6PHIC_2S_3_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L6PHIC_2S_4_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L6PHIC_2S_4_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L6PHIC_2S_4_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L6PHIC_2S_4_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L6PHIC_2S_4_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L6PHIC_neg2S_3_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L6PHIC_neg2S_3_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L6PHIC_neg2S_3_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_L6PHIC_neg2S_3_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L6PHIC_neg2S_3_A_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_L6PHIC_neg2S_3_B_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_L6PHIC_neg2S_3_B_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_L6PHIC_neg2S_3_B_V_dout,
      inputStubs_4_nentries_0_V               => IL_L6PHIC_neg2S_3_B_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_L6PHIC_neg2S_3_B_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_L6PHIC_neg2S_4_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_L6PHIC_neg2S_4_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_L6PHIC_neg2S_4_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_L6PHIC_neg2S_4_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_L6PHIC_neg2S_4_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHICn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L6PHIC_B_L5C_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L6PHIC_B_L5C_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L6PHIC_B_L5C_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L6PHICn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L6PHICn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L6PHICn1_din
  );

  LATCH_VMR_L6PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_L6PHID_bx,
      start => VMR_L6PHID_start
  );

  VMR_L6PHID : entity work.VMR_L6PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_L6PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_L6PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_L6PHID_2S_3_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_L6PHID_2S_3_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_L6PHID_2S_3_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_L6PHID_2S_3_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_L6PHID_2S_3_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_L6PHID_2S_4_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_L6PHID_2S_4_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_L6PHID_2S_4_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_L6PHID_2S_4_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_L6PHID_2S_4_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_L6PHID_neg2S_3_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_L6PHID_neg2S_3_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_L6PHID_neg2S_3_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_L6PHID_neg2S_3_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_L6PHID_neg2S_3_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_L6PHID_neg2S_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_L6PHID_neg2S_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_L6PHID_neg2S_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_L6PHID_neg2S_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_L6PHID_neg2S_4_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_L6PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_L6PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_L6PHIDn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_L6PHID_B_L5D_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_L6PHID_B_L5D_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_L6PHID_B_L5D_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_L6PHIDn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_L6PHIDn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_L6PHIDn1_din
  );

  LATCH_VMR_D1PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D1PHIA_bx,
      start => VMR_D1PHIA_start
  );

  VMR_D1PHIA : entity work.VMR_D1PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D1PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D1PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D1PHIA_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D1PHIA_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D1PHIA_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D1PHIA_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D1PHIA_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D1PHIA_PS10G_4_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D1PHIA_PS10G_4_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D1PHIA_PS10G_4_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_D1PHIA_PS10G_4_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D1PHIA_PS10G_4_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D1PHIA_negPS10G_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D1PHIA_negPS10G_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D1PHIA_negPS10G_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D1PHIA_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D1PHIA_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D1PHIA_negPS10G_4_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D1PHIA_negPS10G_4_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D1PHIA_negPS10G_4_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_D1PHIA_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D1PHIA_negPS10G_4_A_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D1PHIA_2S_5_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D1PHIA_2S_5_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D1PHIA_2S_5_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D1PHIA_2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D1PHIA_2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D1PHIA_neg2S_5_A_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D1PHIA_neg2S_5_A_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D1PHIA_neg2S_5_A_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D1PHIA_neg2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D1PHIA_neg2S_5_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHIAn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D1PHIA_O_L1A_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D1PHIA_O_L1A_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D1PHIA_O_L1A_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_D1PHIA_O_L1B_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_D1PHIA_O_L1B_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_D1PHIA_O_L1B_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_D1PHIA_O_L2A_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_D1PHIA_O_L2A_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_D1PHIA_O_L2A_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D1PHIA_DM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D1PHIA_DM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D1PHIA_DM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D1PHIXn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D1PHIXn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D1PHIXn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_D1PHIXn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_D1PHIXn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_D1PHIXn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_D1PHIXn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_D1PHIXn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_D1PHIXn3_din
  );

  LATCH_VMR_D1PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D1PHIB_bx,
      start => VMR_D1PHIB_start
  );

  VMR_D1PHIB : entity work.VMR_D1PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D1PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D1PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D1PHIB_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D1PHIB_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D1PHIB_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D1PHIB_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D1PHIB_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D1PHIB_PS10G_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D1PHIB_PS10G_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D1PHIB_PS10G_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D1PHIB_PS10G_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D1PHIB_PS10G_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D1PHIB_PS10G_4_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D1PHIB_PS10G_4_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D1PHIB_PS10G_4_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D1PHIB_PS10G_4_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D1PHIB_PS10G_4_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D1PHIB_PS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D1PHIB_PS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D1PHIB_PS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D1PHIB_PS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D1PHIB_PS10G_4_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D1PHIB_negPS10G_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D1PHIB_negPS10G_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D1PHIB_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D1PHIB_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D1PHIB_negPS10G_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D1PHIB_negPS10G_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D1PHIB_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D1PHIB_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D1PHIB_negPS10G_4_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_4_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D1PHIB_negPS10G_4_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D1PHIB_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D1PHIB_negPS10G_4_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D1PHIB_negPS10G_4_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D1PHIB_negPS10G_4_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D1PHIB_negPS10G_4_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D1PHIB_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D1PHIB_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D1PHIB_2S_5_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D1PHIB_2S_5_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D1PHIB_2S_5_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D1PHIB_2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D1PHIB_2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D1PHIB_2S_5_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D1PHIB_2S_5_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D1PHIB_2S_5_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D1PHIB_2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D1PHIB_2S_5_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D1PHIB_neg2S_5_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D1PHIB_neg2S_5_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D1PHIB_neg2S_5_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D1PHIB_neg2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D1PHIB_neg2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D1PHIB_neg2S_5_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D1PHIB_neg2S_5_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D1PHIB_neg2S_5_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D1PHIB_neg2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D1PHIB_neg2S_5_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHIBn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D1PHIB_O_L1C_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D1PHIB_O_L1C_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D1PHIB_O_L1C_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_D1PHIB_O_L1D_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_D1PHIB_O_L1D_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_D1PHIB_O_L1D_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_D1PHIB_O_L2B_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_D1PHIB_O_L2B_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_D1PHIB_O_L2B_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D1PHIB_DM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D1PHIB_DM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D1PHIB_DM_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_D1PHIB_DR_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_D1PHIB_DR_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_D1PHIB_DR_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D1PHIYn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D1PHIYn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D1PHIYn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_D1PHIYn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_D1PHIYn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_D1PHIYn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_D1PHIYn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_D1PHIYn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_D1PHIYn3_din
  );

  LATCH_VMR_D1PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D1PHIC_bx,
      start => VMR_D1PHIC_start
  );

  VMR_D1PHIC : entity work.VMR_D1PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D1PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D1PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D1PHIC_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D1PHIC_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D1PHIC_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D1PHIC_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D1PHIC_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D1PHIC_PS10G_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D1PHIC_PS10G_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D1PHIC_PS10G_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D1PHIC_PS10G_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D1PHIC_PS10G_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D1PHIC_PS10G_4_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D1PHIC_PS10G_4_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D1PHIC_PS10G_4_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D1PHIC_PS10G_4_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D1PHIC_PS10G_4_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D1PHIC_PS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D1PHIC_PS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D1PHIC_PS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D1PHIC_PS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D1PHIC_PS10G_4_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D1PHIC_negPS10G_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D1PHIC_negPS10G_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D1PHIC_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D1PHIC_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D1PHIC_negPS10G_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D1PHIC_negPS10G_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D1PHIC_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D1PHIC_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D1PHIC_negPS10G_4_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_4_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D1PHIC_negPS10G_4_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D1PHIC_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D1PHIC_negPS10G_4_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D1PHIC_negPS10G_4_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D1PHIC_negPS10G_4_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D1PHIC_negPS10G_4_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D1PHIC_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D1PHIC_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D1PHIC_2S_5_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D1PHIC_2S_5_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D1PHIC_2S_5_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D1PHIC_2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D1PHIC_2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D1PHIC_2S_5_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D1PHIC_2S_5_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D1PHIC_2S_5_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D1PHIC_2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D1PHIC_2S_5_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D1PHIC_neg2S_5_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D1PHIC_neg2S_5_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D1PHIC_neg2S_5_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D1PHIC_neg2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D1PHIC_neg2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D1PHIC_neg2S_5_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D1PHIC_neg2S_5_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D1PHIC_neg2S_5_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D1PHIC_neg2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D1PHIC_neg2S_5_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHICn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D1PHIC_O_L1E_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D1PHIC_O_L1E_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D1PHIC_O_L1E_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_D1PHIC_O_L1F_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_D1PHIC_O_L1F_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_D1PHIC_O_L1F_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_D1PHIC_O_L2C_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_D1PHIC_O_L2C_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_D1PHIC_O_L2C_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D1PHIC_DL_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D1PHIC_DL_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D1PHIC_DL_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_D1PHIC_DM_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_D1PHIC_DM_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_D1PHIC_DM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D1PHIZn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D1PHIZn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D1PHIZn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_D1PHIZn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_D1PHIZn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_D1PHIZn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_D1PHIZn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_D1PHIZn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_D1PHIZn3_din
  );

  LATCH_VMR_D1PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D1PHID_bx,
      start => VMR_D1PHID_start
  );

  VMR_D1PHID : entity work.VMR_D1PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D1PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D1PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D1PHID_PS10G_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D1PHID_PS10G_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D1PHID_PS10G_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_D1PHID_PS10G_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D1PHID_PS10G_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D1PHID_PS10G_4_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D1PHID_PS10G_4_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D1PHID_PS10G_4_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D1PHID_PS10G_4_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D1PHID_PS10G_4_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D1PHID_negPS10G_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D1PHID_negPS10G_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D1PHID_negPS10G_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_D1PHID_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D1PHID_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D1PHID_negPS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D1PHID_negPS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D1PHID_negPS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D1PHID_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D1PHID_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D1PHID_2S_5_B_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D1PHID_2S_5_B_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D1PHID_2S_5_B_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D1PHID_2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D1PHID_2S_5_B_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D1PHID_neg2S_5_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D1PHID_neg2S_5_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D1PHID_neg2S_5_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D1PHID_neg2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D1PHID_neg2S_5_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D1PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D1PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D1PHIDn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D1PHID_O_L1G_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D1PHID_O_L1G_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D1PHID_O_L1G_din,
      memoriesAS_2_dataarray_data_V_ce0       => open,
      memoriesAS_2_dataarray_data_V_we0       => AS_D1PHID_O_L1H_wea,
      memoriesAS_2_dataarray_data_V_address0  => AS_D1PHID_O_L1H_writeaddr,
      memoriesAS_2_dataarray_data_V_d0        => AS_D1PHID_O_L1H_din,
      memoriesAS_3_dataarray_data_V_ce0       => open,
      memoriesAS_3_dataarray_data_V_we0       => AS_D1PHID_O_L2D_wea,
      memoriesAS_3_dataarray_data_V_address0  => AS_D1PHID_O_L2D_writeaddr,
      memoriesAS_3_dataarray_data_V_d0        => AS_D1PHID_O_L2D_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D1PHID_DM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D1PHID_DM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D1PHID_DM_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D1PHIWn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D1PHIWn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D1PHIWn1_din,
      memoriesTEO_1_dataarray_0_data_V_ce0       => open,
      memoriesTEO_1_dataarray_0_data_V_we0       => VMSTE_D1PHIWn2_wea,
      memoriesTEO_1_dataarray_0_data_V_address0  => VMSTE_D1PHIWn2_writeaddr,
      memoriesTEO_1_dataarray_0_data_V_d0        => VMSTE_D1PHIWn2_din,
      memoriesTEO_2_dataarray_0_data_V_ce0       => open,
      memoriesTEO_2_dataarray_0_data_V_we0       => VMSTE_D1PHIWn3_wea,
      memoriesTEO_2_dataarray_0_data_V_address0  => VMSTE_D1PHIWn3_writeaddr,
      memoriesTEO_2_dataarray_0_data_V_d0        => VMSTE_D1PHIWn3_din
  );

  LATCH_VMR_D2PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D2PHIA_bx,
      start => VMR_D2PHIA_start
  );

  VMR_D2PHIA : entity work.VMR_D2PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D2PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D2PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D2PHIA_PS10G_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D2PHIA_PS10G_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D2PHIA_PS10G_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D2PHIA_PS10G_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D2PHIA_PS10G_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D2PHIA_PS10G_3_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D2PHIA_PS10G_3_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D2PHIA_PS10G_3_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_D2PHIA_PS10G_3_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D2PHIA_PS10G_3_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D2PHIA_PS_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D2PHIA_PS_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D2PHIA_PS_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D2PHIA_PS_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D2PHIA_PS_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D2PHIA_negPS10G_2_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D2PHIA_negPS10G_2_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D2PHIA_negPS10G_2_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_D2PHIA_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D2PHIA_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D2PHIA_negPS10G_3_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D2PHIA_negPS10G_3_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D2PHIA_negPS10G_3_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D2PHIA_negPS10G_3_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D2PHIA_negPS10G_3_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D2PHIA_negPS_1_A_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D2PHIA_negPS_1_A_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D2PHIA_negPS_1_A_V_dout,
      inputStubs_5_nentries_0_V               => IL_D2PHIA_negPS_1_A_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D2PHIA_negPS_1_A_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D2PHIA_2S_6_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D2PHIA_2S_6_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D2PHIA_2S_6_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D2PHIA_2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D2PHIA_2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D2PHIA_neg2S_6_A_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D2PHIA_neg2S_6_A_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D2PHIA_neg2S_6_A_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D2PHIA_neg2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D2PHIA_neg2S_6_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHIAn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D2PHIA_D_D1A_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D2PHIA_D_D1A_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D2PHIA_D_D1A_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D2PHIAn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D2PHIAn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D2PHIAn1_din
  );

  LATCH_VMR_D2PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D2PHIB_bx,
      start => VMR_D2PHIB_start
  );

  VMR_D2PHIB : entity work.VMR_D2PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D2PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D2PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D2PHIB_PS10G_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D2PHIB_PS10G_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D2PHIB_PS10G_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D2PHIB_PS10G_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D2PHIB_PS10G_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D2PHIB_PS10G_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D2PHIB_PS10G_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D2PHIB_PS10G_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D2PHIB_PS10G_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D2PHIB_PS10G_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D2PHIB_PS10G_3_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D2PHIB_PS10G_3_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D2PHIB_PS10G_3_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D2PHIB_PS10G_3_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D2PHIB_PS10G_3_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D2PHIB_PS10G_3_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D2PHIB_PS10G_3_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D2PHIB_PS10G_3_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D2PHIB_PS10G_3_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D2PHIB_PS10G_3_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D2PHIB_PS_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D2PHIB_PS_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D2PHIB_PS_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D2PHIB_PS_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D2PHIB_PS_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D2PHIB_PS_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D2PHIB_PS_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D2PHIB_PS_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D2PHIB_PS_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D2PHIB_PS_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D2PHIB_negPS10G_2_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_2_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D2PHIB_negPS10G_2_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D2PHIB_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D2PHIB_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D2PHIB_negPS10G_2_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_2_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D2PHIB_negPS10G_2_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D2PHIB_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D2PHIB_negPS10G_2_B_AV_dout_nent(1),
      inputStubs_8_dataarray_data_V_ce0       => IL_D2PHIB_negPS10G_3_A_enb,
      inputStubs_8_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_3_A_V_readaddr,
      inputStubs_8_dataarray_data_V_q0        => IL_D2PHIB_negPS10G_3_A_V_dout,
      inputStubs_8_nentries_0_V               => IL_D2PHIB_negPS10G_3_A_AV_dout_nent(0),
      inputStubs_8_nentries_1_V               => IL_D2PHIB_negPS10G_3_A_AV_dout_nent(1),
      inputStubs_9_dataarray_data_V_ce0       => IL_D2PHIB_negPS10G_3_B_enb,
      inputStubs_9_dataarray_data_V_address0  => IL_D2PHIB_negPS10G_3_B_V_readaddr,
      inputStubs_9_dataarray_data_V_q0        => IL_D2PHIB_negPS10G_3_B_V_dout,
      inputStubs_9_nentries_0_V               => IL_D2PHIB_negPS10G_3_B_AV_dout_nent(0),
      inputStubs_9_nentries_1_V               => IL_D2PHIB_negPS10G_3_B_AV_dout_nent(1),
      inputStubs_10_dataarray_data_V_ce0       => IL_D2PHIB_negPS_1_A_enb,
      inputStubs_10_dataarray_data_V_address0  => IL_D2PHIB_negPS_1_A_V_readaddr,
      inputStubs_10_dataarray_data_V_q0        => IL_D2PHIB_negPS_1_A_V_dout,
      inputStubs_10_nentries_0_V               => IL_D2PHIB_negPS_1_A_AV_dout_nent(0),
      inputStubs_10_nentries_1_V               => IL_D2PHIB_negPS_1_A_AV_dout_nent(1),
      inputStubs_11_dataarray_data_V_ce0       => IL_D2PHIB_negPS_1_B_enb,
      inputStubs_11_dataarray_data_V_address0  => IL_D2PHIB_negPS_1_B_V_readaddr,
      inputStubs_11_dataarray_data_V_q0        => IL_D2PHIB_negPS_1_B_V_dout,
      inputStubs_11_nentries_0_V               => IL_D2PHIB_negPS_1_B_AV_dout_nent(0),
      inputStubs_11_nentries_1_V               => IL_D2PHIB_negPS_1_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D2PHIB_2S_6_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D2PHIB_2S_6_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D2PHIB_2S_6_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D2PHIB_2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D2PHIB_2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D2PHIB_2S_6_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D2PHIB_2S_6_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D2PHIB_2S_6_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D2PHIB_2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D2PHIB_2S_6_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D2PHIB_neg2S_6_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D2PHIB_neg2S_6_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D2PHIB_neg2S_6_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D2PHIB_neg2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D2PHIB_neg2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D2PHIB_neg2S_6_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D2PHIB_neg2S_6_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D2PHIB_neg2S_6_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D2PHIB_neg2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D2PHIB_neg2S_6_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHIBn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D2PHIB_D_D1B_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D2PHIB_D_D1B_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D2PHIB_D_D1B_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D2PHIBn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D2PHIBn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D2PHIBn1_din
  );

  LATCH_VMR_D2PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D2PHIC_bx,
      start => VMR_D2PHIC_start
  );

  VMR_D2PHIC : entity work.VMR_D2PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D2PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D2PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D2PHIC_PS10G_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D2PHIC_PS10G_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D2PHIC_PS10G_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D2PHIC_PS10G_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D2PHIC_PS10G_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D2PHIC_PS10G_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D2PHIC_PS10G_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D2PHIC_PS10G_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D2PHIC_PS10G_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D2PHIC_PS10G_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D2PHIC_PS10G_3_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D2PHIC_PS10G_3_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D2PHIC_PS10G_3_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D2PHIC_PS10G_3_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D2PHIC_PS10G_3_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D2PHIC_PS10G_3_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D2PHIC_PS10G_3_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D2PHIC_PS10G_3_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D2PHIC_PS10G_3_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D2PHIC_PS10G_3_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D2PHIC_PS_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D2PHIC_PS_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D2PHIC_PS_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D2PHIC_PS_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D2PHIC_PS_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D2PHIC_PS_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D2PHIC_PS_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D2PHIC_PS_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D2PHIC_PS_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D2PHIC_PS_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D2PHIC_negPS10G_2_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_2_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D2PHIC_negPS10G_2_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D2PHIC_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D2PHIC_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D2PHIC_negPS10G_2_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_2_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D2PHIC_negPS10G_2_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D2PHIC_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D2PHIC_negPS10G_2_B_AV_dout_nent(1),
      inputStubs_8_dataarray_data_V_ce0       => IL_D2PHIC_negPS10G_3_A_enb,
      inputStubs_8_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_3_A_V_readaddr,
      inputStubs_8_dataarray_data_V_q0        => IL_D2PHIC_negPS10G_3_A_V_dout,
      inputStubs_8_nentries_0_V               => IL_D2PHIC_negPS10G_3_A_AV_dout_nent(0),
      inputStubs_8_nentries_1_V               => IL_D2PHIC_negPS10G_3_A_AV_dout_nent(1),
      inputStubs_9_dataarray_data_V_ce0       => IL_D2PHIC_negPS10G_3_B_enb,
      inputStubs_9_dataarray_data_V_address0  => IL_D2PHIC_negPS10G_3_B_V_readaddr,
      inputStubs_9_dataarray_data_V_q0        => IL_D2PHIC_negPS10G_3_B_V_dout,
      inputStubs_9_nentries_0_V               => IL_D2PHIC_negPS10G_3_B_AV_dout_nent(0),
      inputStubs_9_nentries_1_V               => IL_D2PHIC_negPS10G_3_B_AV_dout_nent(1),
      inputStubs_10_dataarray_data_V_ce0       => IL_D2PHIC_negPS_1_A_enb,
      inputStubs_10_dataarray_data_V_address0  => IL_D2PHIC_negPS_1_A_V_readaddr,
      inputStubs_10_dataarray_data_V_q0        => IL_D2PHIC_negPS_1_A_V_dout,
      inputStubs_10_nentries_0_V               => IL_D2PHIC_negPS_1_A_AV_dout_nent(0),
      inputStubs_10_nentries_1_V               => IL_D2PHIC_negPS_1_A_AV_dout_nent(1),
      inputStubs_11_dataarray_data_V_ce0       => IL_D2PHIC_negPS_1_B_enb,
      inputStubs_11_dataarray_data_V_address0  => IL_D2PHIC_negPS_1_B_V_readaddr,
      inputStubs_11_dataarray_data_V_q0        => IL_D2PHIC_negPS_1_B_V_dout,
      inputStubs_11_nentries_0_V               => IL_D2PHIC_negPS_1_B_AV_dout_nent(0),
      inputStubs_11_nentries_1_V               => IL_D2PHIC_negPS_1_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D2PHIC_2S_6_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D2PHIC_2S_6_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D2PHIC_2S_6_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D2PHIC_2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D2PHIC_2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D2PHIC_2S_6_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D2PHIC_2S_6_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D2PHIC_2S_6_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D2PHIC_2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D2PHIC_2S_6_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D2PHIC_neg2S_6_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D2PHIC_neg2S_6_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D2PHIC_neg2S_6_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D2PHIC_neg2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D2PHIC_neg2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D2PHIC_neg2S_6_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D2PHIC_neg2S_6_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D2PHIC_neg2S_6_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D2PHIC_neg2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D2PHIC_neg2S_6_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHICn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D2PHIC_D_D1C_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D2PHIC_D_D1C_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D2PHIC_D_D1C_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D2PHICn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D2PHICn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D2PHICn1_din
  );

  LATCH_VMR_D2PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D2PHID_bx,
      start => VMR_D2PHID_start
  );

  VMR_D2PHID : entity work.VMR_D2PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D2PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D2PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D2PHID_PS10G_2_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D2PHID_PS10G_2_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D2PHID_PS10G_2_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_D2PHID_PS10G_2_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D2PHID_PS10G_2_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D2PHID_PS10G_3_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D2PHID_PS10G_3_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D2PHID_PS10G_3_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D2PHID_PS10G_3_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D2PHID_PS10G_3_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D2PHID_PS_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D2PHID_PS_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D2PHID_PS_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_D2PHID_PS_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D2PHID_PS_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D2PHID_negPS10G_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D2PHID_negPS10G_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D2PHID_negPS10G_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D2PHID_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D2PHID_negPS10G_2_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D2PHID_negPS10G_3_B_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D2PHID_negPS10G_3_B_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D2PHID_negPS10G_3_B_V_dout,
      inputStubs_4_nentries_0_V               => IL_D2PHID_negPS10G_3_B_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D2PHID_negPS10G_3_B_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D2PHID_negPS_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D2PHID_negPS_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D2PHID_negPS_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D2PHID_negPS_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D2PHID_negPS_1_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D2PHID_2S_6_B_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D2PHID_2S_6_B_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D2PHID_2S_6_B_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D2PHID_2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D2PHID_2S_6_B_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D2PHID_neg2S_6_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D2PHID_neg2S_6_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D2PHID_neg2S_6_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D2PHID_neg2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D2PHID_neg2S_6_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D2PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D2PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D2PHIDn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D2PHID_D_D1D_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D2PHID_D_D1D_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D2PHID_D_D1D_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D2PHIDn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D2PHIDn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D2PHIDn1_din
  );

  LATCH_VMR_D3PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D3PHIA_bx,
      start => VMR_D3PHIA_start
  );

  VMR_D3PHIA : entity work.VMR_D3PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D3PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D3PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D3PHIA_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D3PHIA_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D3PHIA_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D3PHIA_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D3PHIA_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D3PHIA_PS10G_4_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D3PHIA_PS10G_4_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D3PHIA_PS10G_4_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_D3PHIA_PS10G_4_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D3PHIA_PS10G_4_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D3PHIA_negPS10G_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D3PHIA_negPS10G_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D3PHIA_negPS10G_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D3PHIA_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D3PHIA_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D3PHIA_negPS10G_4_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D3PHIA_negPS10G_4_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D3PHIA_negPS10G_4_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_D3PHIA_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D3PHIA_negPS10G_4_A_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D3PHIA_2S_4_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D3PHIA_2S_4_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D3PHIA_2S_4_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D3PHIA_2S_4_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D3PHIA_2S_4_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D3PHIA_neg2S_4_A_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D3PHIA_neg2S_4_A_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D3PHIA_neg2S_4_A_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D3PHIA_neg2S_4_A_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D3PHIA_neg2S_4_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHIAn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D3PHIA_DM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D3PHIA_DM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D3PHIA_DM_din
  );

  LATCH_VMR_D3PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D3PHIB_bx,
      start => VMR_D3PHIB_start
  );

  VMR_D3PHIB : entity work.VMR_D3PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D3PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D3PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D3PHIB_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D3PHIB_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D3PHIB_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D3PHIB_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D3PHIB_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D3PHIB_PS10G_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D3PHIB_PS10G_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D3PHIB_PS10G_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D3PHIB_PS10G_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D3PHIB_PS10G_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D3PHIB_PS10G_4_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D3PHIB_PS10G_4_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D3PHIB_PS10G_4_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D3PHIB_PS10G_4_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D3PHIB_PS10G_4_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D3PHIB_PS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D3PHIB_PS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D3PHIB_PS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D3PHIB_PS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D3PHIB_PS10G_4_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D3PHIB_negPS10G_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D3PHIB_negPS10G_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D3PHIB_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D3PHIB_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D3PHIB_negPS10G_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D3PHIB_negPS10G_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D3PHIB_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D3PHIB_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D3PHIB_negPS10G_4_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_4_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D3PHIB_negPS10G_4_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D3PHIB_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D3PHIB_negPS10G_4_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D3PHIB_negPS10G_4_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D3PHIB_negPS10G_4_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D3PHIB_negPS10G_4_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D3PHIB_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D3PHIB_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D3PHIB_2S_4_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D3PHIB_2S_4_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D3PHIB_2S_4_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D3PHIB_2S_4_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D3PHIB_2S_4_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D3PHIB_2S_4_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D3PHIB_2S_4_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D3PHIB_2S_4_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D3PHIB_2S_4_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D3PHIB_2S_4_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D3PHIB_neg2S_4_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D3PHIB_neg2S_4_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D3PHIB_neg2S_4_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D3PHIB_neg2S_4_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D3PHIB_neg2S_4_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D3PHIB_neg2S_4_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D3PHIB_neg2S_4_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D3PHIB_neg2S_4_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D3PHIB_neg2S_4_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D3PHIB_neg2S_4_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHIBn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D3PHIB_DM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D3PHIB_DM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D3PHIB_DM_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_D3PHIB_DR_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_D3PHIB_DR_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_D3PHIB_DR_din
  );

  LATCH_VMR_D3PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D3PHIC_bx,
      start => VMR_D3PHIC_start
  );

  VMR_D3PHIC : entity work.VMR_D3PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D3PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D3PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D3PHIC_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D3PHIC_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D3PHIC_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D3PHIC_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D3PHIC_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D3PHIC_PS10G_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D3PHIC_PS10G_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D3PHIC_PS10G_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D3PHIC_PS10G_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D3PHIC_PS10G_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D3PHIC_PS10G_4_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D3PHIC_PS10G_4_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D3PHIC_PS10G_4_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D3PHIC_PS10G_4_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D3PHIC_PS10G_4_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D3PHIC_PS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D3PHIC_PS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D3PHIC_PS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D3PHIC_PS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D3PHIC_PS10G_4_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D3PHIC_negPS10G_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D3PHIC_negPS10G_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D3PHIC_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D3PHIC_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D3PHIC_negPS10G_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D3PHIC_negPS10G_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D3PHIC_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D3PHIC_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D3PHIC_negPS10G_4_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_4_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D3PHIC_negPS10G_4_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D3PHIC_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D3PHIC_negPS10G_4_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D3PHIC_negPS10G_4_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D3PHIC_negPS10G_4_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D3PHIC_negPS10G_4_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D3PHIC_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D3PHIC_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D3PHIC_2S_4_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D3PHIC_2S_4_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D3PHIC_2S_4_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D3PHIC_2S_4_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D3PHIC_2S_4_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D3PHIC_2S_4_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D3PHIC_2S_4_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D3PHIC_2S_4_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D3PHIC_2S_4_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D3PHIC_2S_4_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D3PHIC_neg2S_4_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D3PHIC_neg2S_4_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D3PHIC_neg2S_4_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D3PHIC_neg2S_4_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D3PHIC_neg2S_4_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D3PHIC_neg2S_4_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D3PHIC_neg2S_4_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D3PHIC_neg2S_4_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D3PHIC_neg2S_4_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D3PHIC_neg2S_4_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHICn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D3PHIC_DL_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D3PHIC_DL_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D3PHIC_DL_din,
      memoriesASInner_1_dataarray_data_V_ce0       => open,
      memoriesASInner_1_dataarray_data_V_we0       => AS_D3PHIC_DM_wea,
      memoriesASInner_1_dataarray_data_V_address0  => AS_D3PHIC_DM_writeaddr,
      memoriesASInner_1_dataarray_data_V_d0        => AS_D3PHIC_DM_din
  );

  LATCH_VMR_D3PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D3PHID_bx,
      start => VMR_D3PHID_start
  );

  VMR_D3PHID : entity work.VMR_D3PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D3PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D3PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D3PHID_PS10G_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D3PHID_PS10G_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D3PHID_PS10G_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_D3PHID_PS10G_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D3PHID_PS10G_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D3PHID_PS10G_4_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D3PHID_PS10G_4_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D3PHID_PS10G_4_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D3PHID_PS10G_4_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D3PHID_PS10G_4_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D3PHID_negPS10G_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D3PHID_negPS10G_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D3PHID_negPS10G_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_D3PHID_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D3PHID_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D3PHID_negPS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D3PHID_negPS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D3PHID_negPS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D3PHID_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D3PHID_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D3PHID_2S_4_B_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D3PHID_2S_4_B_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D3PHID_2S_4_B_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D3PHID_2S_4_B_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D3PHID_2S_4_B_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D3PHID_neg2S_4_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D3PHID_neg2S_4_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D3PHID_neg2S_4_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D3PHID_neg2S_4_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D3PHID_neg2S_4_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D3PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D3PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D3PHIDn1_din,
      memoriesASInner_0_dataarray_data_V_ce0       => open,
      memoriesASInner_0_dataarray_data_V_we0       => AS_D3PHID_DM_wea,
      memoriesASInner_0_dataarray_data_V_address0  => AS_D3PHID_DM_writeaddr,
      memoriesASInner_0_dataarray_data_V_d0        => AS_D3PHID_DM_din
  );

  LATCH_VMR_D4PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D4PHIA_bx,
      start => VMR_D4PHIA_start
  );

  VMR_D4PHIA : entity work.VMR_D4PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D4PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D4PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D4PHIA_PS10G_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D4PHIA_PS10G_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D4PHIA_PS10G_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D4PHIA_PS10G_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D4PHIA_PS10G_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D4PHIA_PS_2_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D4PHIA_PS_2_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D4PHIA_PS_2_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_D4PHIA_PS_2_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D4PHIA_PS_2_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D4PHIA_negPS10G_2_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D4PHIA_negPS10G_2_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D4PHIA_negPS10G_2_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D4PHIA_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D4PHIA_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D4PHIA_negPS_2_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D4PHIA_negPS_2_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D4PHIA_negPS_2_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_D4PHIA_negPS_2_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D4PHIA_negPS_2_A_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D4PHIA_2S_5_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D4PHIA_2S_5_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D4PHIA_2S_5_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D4PHIA_2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D4PHIA_2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D4PHIA_neg2S_5_A_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D4PHIA_neg2S_5_A_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D4PHIA_neg2S_5_A_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D4PHIA_neg2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D4PHIA_neg2S_5_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHIAn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D4PHIA_D_D3A_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D4PHIA_D_D3A_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D4PHIA_D_D3A_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D4PHIAn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D4PHIAn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D4PHIAn1_din
  );

  LATCH_VMR_D4PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D4PHIB_bx,
      start => VMR_D4PHIB_start
  );

  VMR_D4PHIB : entity work.VMR_D4PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D4PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D4PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D4PHIB_PS10G_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D4PHIB_PS10G_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D4PHIB_PS10G_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D4PHIB_PS10G_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D4PHIB_PS10G_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D4PHIB_PS10G_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D4PHIB_PS10G_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D4PHIB_PS10G_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D4PHIB_PS10G_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D4PHIB_PS10G_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D4PHIB_PS_2_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D4PHIB_PS_2_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D4PHIB_PS_2_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D4PHIB_PS_2_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D4PHIB_PS_2_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D4PHIB_PS_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D4PHIB_PS_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D4PHIB_PS_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D4PHIB_PS_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D4PHIB_PS_2_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D4PHIB_negPS10G_2_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D4PHIB_negPS10G_2_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D4PHIB_negPS10G_2_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D4PHIB_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D4PHIB_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D4PHIB_negPS10G_2_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D4PHIB_negPS10G_2_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D4PHIB_negPS10G_2_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D4PHIB_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D4PHIB_negPS10G_2_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D4PHIB_negPS_2_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D4PHIB_negPS_2_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D4PHIB_negPS_2_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D4PHIB_negPS_2_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D4PHIB_negPS_2_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D4PHIB_negPS_2_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D4PHIB_negPS_2_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D4PHIB_negPS_2_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D4PHIB_negPS_2_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D4PHIB_negPS_2_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D4PHIB_2S_5_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D4PHIB_2S_5_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D4PHIB_2S_5_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D4PHIB_2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D4PHIB_2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D4PHIB_2S_5_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D4PHIB_2S_5_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D4PHIB_2S_5_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D4PHIB_2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D4PHIB_2S_5_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D4PHIB_neg2S_5_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D4PHIB_neg2S_5_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D4PHIB_neg2S_5_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D4PHIB_neg2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D4PHIB_neg2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D4PHIB_neg2S_5_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D4PHIB_neg2S_5_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D4PHIB_neg2S_5_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D4PHIB_neg2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D4PHIB_neg2S_5_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHIBn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D4PHIB_D_D3B_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D4PHIB_D_D3B_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D4PHIB_D_D3B_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D4PHIBn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D4PHIBn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D4PHIBn1_din
  );

  LATCH_VMR_D4PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D4PHIC_bx,
      start => VMR_D4PHIC_start
  );

  VMR_D4PHIC : entity work.VMR_D4PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D4PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D4PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D4PHIC_PS10G_2_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D4PHIC_PS10G_2_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D4PHIC_PS10G_2_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D4PHIC_PS10G_2_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D4PHIC_PS10G_2_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D4PHIC_PS10G_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D4PHIC_PS10G_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D4PHIC_PS10G_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D4PHIC_PS10G_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D4PHIC_PS10G_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D4PHIC_PS_2_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D4PHIC_PS_2_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D4PHIC_PS_2_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D4PHIC_PS_2_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D4PHIC_PS_2_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D4PHIC_PS_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D4PHIC_PS_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D4PHIC_PS_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D4PHIC_PS_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D4PHIC_PS_2_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D4PHIC_negPS10G_2_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D4PHIC_negPS10G_2_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D4PHIC_negPS10G_2_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D4PHIC_negPS10G_2_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D4PHIC_negPS10G_2_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D4PHIC_negPS10G_2_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D4PHIC_negPS10G_2_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D4PHIC_negPS10G_2_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D4PHIC_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D4PHIC_negPS10G_2_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D4PHIC_negPS_2_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D4PHIC_negPS_2_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D4PHIC_negPS_2_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D4PHIC_negPS_2_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D4PHIC_negPS_2_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D4PHIC_negPS_2_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D4PHIC_negPS_2_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D4PHIC_negPS_2_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D4PHIC_negPS_2_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D4PHIC_negPS_2_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D4PHIC_2S_5_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D4PHIC_2S_5_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D4PHIC_2S_5_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D4PHIC_2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D4PHIC_2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D4PHIC_2S_5_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D4PHIC_2S_5_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D4PHIC_2S_5_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D4PHIC_2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D4PHIC_2S_5_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D4PHIC_neg2S_5_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D4PHIC_neg2S_5_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D4PHIC_neg2S_5_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D4PHIC_neg2S_5_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D4PHIC_neg2S_5_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D4PHIC_neg2S_5_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D4PHIC_neg2S_5_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D4PHIC_neg2S_5_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D4PHIC_neg2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D4PHIC_neg2S_5_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHICn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D4PHIC_D_D3C_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D4PHIC_D_D3C_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D4PHIC_D_D3C_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D4PHICn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D4PHICn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D4PHICn1_din
  );

  LATCH_VMR_D4PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D4PHID_bx,
      start => VMR_D4PHID_start
  );

  VMR_D4PHID : entity work.VMR_D4PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D4PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D4PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D4PHID_PS10G_2_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D4PHID_PS10G_2_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D4PHID_PS10G_2_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_D4PHID_PS10G_2_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D4PHID_PS10G_2_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D4PHID_PS_2_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D4PHID_PS_2_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D4PHID_PS_2_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D4PHID_PS_2_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D4PHID_PS_2_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D4PHID_negPS10G_2_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D4PHID_negPS10G_2_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D4PHID_negPS10G_2_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_D4PHID_negPS10G_2_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D4PHID_negPS10G_2_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D4PHID_negPS_2_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D4PHID_negPS_2_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D4PHID_negPS_2_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D4PHID_negPS_2_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D4PHID_negPS_2_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D4PHID_2S_5_B_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D4PHID_2S_5_B_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D4PHID_2S_5_B_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D4PHID_2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D4PHID_2S_5_B_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D4PHID_neg2S_5_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D4PHID_neg2S_5_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D4PHID_neg2S_5_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D4PHID_neg2S_5_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D4PHID_neg2S_5_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D4PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D4PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D4PHIDn1_din,
      memoriesAS_1_dataarray_data_V_ce0       => open,
      memoriesAS_1_dataarray_data_V_we0       => AS_D4PHID_D_D3D_wea,
      memoriesAS_1_dataarray_data_V_address0  => AS_D4PHID_D_D3D_writeaddr,
      memoriesAS_1_dataarray_data_V_d0        => AS_D4PHID_D_D3D_din,
      memoriesTEO_0_dataarray_0_data_V_ce0       => open,
      memoriesTEO_0_dataarray_0_data_V_we0       => VMSTE_D4PHIDn1_wea,
      memoriesTEO_0_dataarray_0_data_V_address0  => VMSTE_D4PHIDn1_writeaddr,
      memoriesTEO_0_dataarray_0_data_V_d0        => VMSTE_D4PHIDn1_din
  );

  LATCH_VMR_D5PHIA: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D5PHIA_bx,
      start => VMR_D5PHIA_start
  );

  VMR_D5PHIA : entity work.VMR_D5PHIA
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D5PHIA_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D5PHIA_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D5PHIA_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D5PHIA_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D5PHIA_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D5PHIA_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D5PHIA_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D5PHIA_PS10G_4_A_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D5PHIA_PS10G_4_A_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D5PHIA_PS10G_4_A_V_dout,
      inputStubs_1_nentries_0_V               => IL_D5PHIA_PS10G_4_A_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D5PHIA_PS10G_4_A_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D5PHIA_negPS10G_1_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D5PHIA_negPS10G_1_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D5PHIA_negPS10G_1_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D5PHIA_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D5PHIA_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D5PHIA_negPS10G_4_A_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D5PHIA_negPS10G_4_A_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D5PHIA_negPS10G_4_A_V_dout,
      inputStubs_3_nentries_0_V               => IL_D5PHIA_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D5PHIA_negPS10G_4_A_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D5PHIA_2S_6_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D5PHIA_2S_6_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D5PHIA_2S_6_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D5PHIA_2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D5PHIA_2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D5PHIA_neg2S_6_A_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D5PHIA_neg2S_6_A_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D5PHIA_neg2S_6_A_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D5PHIA_neg2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D5PHIA_neg2S_6_A_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHIAn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHIAn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHIAn1_din
  );

  LATCH_VMR_D5PHIB: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D5PHIB_bx,
      start => VMR_D5PHIB_start
  );

  VMR_D5PHIB : entity work.VMR_D5PHIB
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D5PHIB_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D5PHIB_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D5PHIB_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D5PHIB_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D5PHIB_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D5PHIB_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D5PHIB_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D5PHIB_PS10G_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D5PHIB_PS10G_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D5PHIB_PS10G_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D5PHIB_PS10G_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D5PHIB_PS10G_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D5PHIB_PS10G_4_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D5PHIB_PS10G_4_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D5PHIB_PS10G_4_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D5PHIB_PS10G_4_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D5PHIB_PS10G_4_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D5PHIB_PS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D5PHIB_PS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D5PHIB_PS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D5PHIB_PS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D5PHIB_PS10G_4_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D5PHIB_negPS10G_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D5PHIB_negPS10G_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D5PHIB_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D5PHIB_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D5PHIB_negPS10G_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D5PHIB_negPS10G_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D5PHIB_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D5PHIB_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D5PHIB_negPS10G_4_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_4_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D5PHIB_negPS10G_4_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D5PHIB_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D5PHIB_negPS10G_4_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D5PHIB_negPS10G_4_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D5PHIB_negPS10G_4_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D5PHIB_negPS10G_4_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D5PHIB_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D5PHIB_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D5PHIB_2S_6_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D5PHIB_2S_6_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D5PHIB_2S_6_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D5PHIB_2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D5PHIB_2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D5PHIB_2S_6_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D5PHIB_2S_6_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D5PHIB_2S_6_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D5PHIB_2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D5PHIB_2S_6_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D5PHIB_neg2S_6_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D5PHIB_neg2S_6_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D5PHIB_neg2S_6_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D5PHIB_neg2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D5PHIB_neg2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D5PHIB_neg2S_6_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D5PHIB_neg2S_6_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D5PHIB_neg2S_6_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D5PHIB_neg2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D5PHIB_neg2S_6_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHIBn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHIBn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHIBn1_din
  );

  LATCH_VMR_D5PHIC: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D5PHIC_bx,
      start => VMR_D5PHIC_start
  );

  VMR_D5PHIC : entity work.VMR_D5PHIC
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D5PHIC_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D5PHIC_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D5PHIC_PS10G_1_A_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D5PHIC_PS10G_1_A_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D5PHIC_PS10G_1_A_V_dout,
      inputStubs_0_nentries_0_V               => IL_D5PHIC_PS10G_1_A_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D5PHIC_PS10G_1_A_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D5PHIC_PS10G_1_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D5PHIC_PS10G_1_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D5PHIC_PS10G_1_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D5PHIC_PS10G_1_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D5PHIC_PS10G_1_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D5PHIC_PS10G_4_A_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D5PHIC_PS10G_4_A_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D5PHIC_PS10G_4_A_V_dout,
      inputStubs_2_nentries_0_V               => IL_D5PHIC_PS10G_4_A_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D5PHIC_PS10G_4_A_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D5PHIC_PS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D5PHIC_PS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D5PHIC_PS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D5PHIC_PS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D5PHIC_PS10G_4_B_AV_dout_nent(1),
      inputStubs_4_dataarray_data_V_ce0       => IL_D5PHIC_negPS10G_1_A_enb,
      inputStubs_4_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_1_A_V_readaddr,
      inputStubs_4_dataarray_data_V_q0        => IL_D5PHIC_negPS10G_1_A_V_dout,
      inputStubs_4_nentries_0_V               => IL_D5PHIC_negPS10G_1_A_AV_dout_nent(0),
      inputStubs_4_nentries_1_V               => IL_D5PHIC_negPS10G_1_A_AV_dout_nent(1),
      inputStubs_5_dataarray_data_V_ce0       => IL_D5PHIC_negPS10G_1_B_enb,
      inputStubs_5_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_1_B_V_readaddr,
      inputStubs_5_dataarray_data_V_q0        => IL_D5PHIC_negPS10G_1_B_V_dout,
      inputStubs_5_nentries_0_V               => IL_D5PHIC_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_5_nentries_1_V               => IL_D5PHIC_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_6_dataarray_data_V_ce0       => IL_D5PHIC_negPS10G_4_A_enb,
      inputStubs_6_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_4_A_V_readaddr,
      inputStubs_6_dataarray_data_V_q0        => IL_D5PHIC_negPS10G_4_A_V_dout,
      inputStubs_6_nentries_0_V               => IL_D5PHIC_negPS10G_4_A_AV_dout_nent(0),
      inputStubs_6_nentries_1_V               => IL_D5PHIC_negPS10G_4_A_AV_dout_nent(1),
      inputStubs_7_dataarray_data_V_ce0       => IL_D5PHIC_negPS10G_4_B_enb,
      inputStubs_7_dataarray_data_V_address0  => IL_D5PHIC_negPS10G_4_B_V_readaddr,
      inputStubs_7_dataarray_data_V_q0        => IL_D5PHIC_negPS10G_4_B_V_dout,
      inputStubs_7_nentries_0_V               => IL_D5PHIC_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_7_nentries_1_V               => IL_D5PHIC_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D5PHIC_2S_6_A_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D5PHIC_2S_6_A_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D5PHIC_2S_6_A_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D5PHIC_2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D5PHIC_2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D5PHIC_2S_6_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D5PHIC_2S_6_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D5PHIC_2S_6_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D5PHIC_2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D5PHIC_2S_6_B_AV_dout_nent(1),
      inputStubsDisk2S_2_dataarray_data_V_ce0       => IL_D5PHIC_neg2S_6_A_enb,
      inputStubsDisk2S_2_dataarray_data_V_address0  => IL_D5PHIC_neg2S_6_A_V_readaddr,
      inputStubsDisk2S_2_dataarray_data_V_q0        => IL_D5PHIC_neg2S_6_A_V_dout,
      inputStubsDisk2S_2_nentries_0_V               => IL_D5PHIC_neg2S_6_A_AV_dout_nent(0),
      inputStubsDisk2S_2_nentries_1_V               => IL_D5PHIC_neg2S_6_A_AV_dout_nent(1),
      inputStubsDisk2S_3_dataarray_data_V_ce0       => IL_D5PHIC_neg2S_6_B_enb,
      inputStubsDisk2S_3_dataarray_data_V_address0  => IL_D5PHIC_neg2S_6_B_V_readaddr,
      inputStubsDisk2S_3_dataarray_data_V_q0        => IL_D5PHIC_neg2S_6_B_V_dout,
      inputStubsDisk2S_3_nentries_0_V               => IL_D5PHIC_neg2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_3_nentries_1_V               => IL_D5PHIC_neg2S_6_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHICn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHICn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHICn1_din
  );

  LATCH_VMR_D5PHID: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => IR_done,
      bx_out => IR_bx_out,
      bx => VMR_D5PHID_bx,
      start => VMR_D5PHID_start
  );

  VMR_D5PHID : entity work.VMR_D5PHID
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => VMR_D5PHID_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => VMR_D5PHID_bx,
      inputStubs_0_dataarray_data_V_ce0       => IL_D5PHID_PS10G_1_B_enb,
      inputStubs_0_dataarray_data_V_address0  => IL_D5PHID_PS10G_1_B_V_readaddr,
      inputStubs_0_dataarray_data_V_q0        => IL_D5PHID_PS10G_1_B_V_dout,
      inputStubs_0_nentries_0_V               => IL_D5PHID_PS10G_1_B_AV_dout_nent(0),
      inputStubs_0_nentries_1_V               => IL_D5PHID_PS10G_1_B_AV_dout_nent(1),
      inputStubs_1_dataarray_data_V_ce0       => IL_D5PHID_PS10G_4_B_enb,
      inputStubs_1_dataarray_data_V_address0  => IL_D5PHID_PS10G_4_B_V_readaddr,
      inputStubs_1_dataarray_data_V_q0        => IL_D5PHID_PS10G_4_B_V_dout,
      inputStubs_1_nentries_0_V               => IL_D5PHID_PS10G_4_B_AV_dout_nent(0),
      inputStubs_1_nentries_1_V               => IL_D5PHID_PS10G_4_B_AV_dout_nent(1),
      inputStubs_2_dataarray_data_V_ce0       => IL_D5PHID_negPS10G_1_B_enb,
      inputStubs_2_dataarray_data_V_address0  => IL_D5PHID_negPS10G_1_B_V_readaddr,
      inputStubs_2_dataarray_data_V_q0        => IL_D5PHID_negPS10G_1_B_V_dout,
      inputStubs_2_nentries_0_V               => IL_D5PHID_negPS10G_1_B_AV_dout_nent(0),
      inputStubs_2_nentries_1_V               => IL_D5PHID_negPS10G_1_B_AV_dout_nent(1),
      inputStubs_3_dataarray_data_V_ce0       => IL_D5PHID_negPS10G_4_B_enb,
      inputStubs_3_dataarray_data_V_address0  => IL_D5PHID_negPS10G_4_B_V_readaddr,
      inputStubs_3_dataarray_data_V_q0        => IL_D5PHID_negPS10G_4_B_V_dout,
      inputStubs_3_nentries_0_V               => IL_D5PHID_negPS10G_4_B_AV_dout_nent(0),
      inputStubs_3_nentries_1_V               => IL_D5PHID_negPS10G_4_B_AV_dout_nent(1),
      inputStubsDisk2S_0_dataarray_data_V_ce0       => IL_D5PHID_2S_6_B_enb,
      inputStubsDisk2S_0_dataarray_data_V_address0  => IL_D5PHID_2S_6_B_V_readaddr,
      inputStubsDisk2S_0_dataarray_data_V_q0        => IL_D5PHID_2S_6_B_V_dout,
      inputStubsDisk2S_0_nentries_0_V               => IL_D5PHID_2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_0_nentries_1_V               => IL_D5PHID_2S_6_B_AV_dout_nent(1),
      inputStubsDisk2S_1_dataarray_data_V_ce0       => IL_D5PHID_neg2S_6_B_enb,
      inputStubsDisk2S_1_dataarray_data_V_address0  => IL_D5PHID_neg2S_6_B_V_readaddr,
      inputStubsDisk2S_1_dataarray_data_V_q0        => IL_D5PHID_neg2S_6_B_V_dout,
      inputStubsDisk2S_1_nentries_0_V               => IL_D5PHID_neg2S_6_B_AV_dout_nent(0),
      inputStubsDisk2S_1_nentries_1_V               => IL_D5PHID_neg2S_6_B_AV_dout_nent(1),
      memoriesAS_0_dataarray_data_V_ce0       => open,
      memoriesAS_0_dataarray_data_V_we0       => AS_D5PHIDn1_wea,
      memoriesAS_0_dataarray_data_V_address0  => AS_D5PHIDn1_writeaddr,
      memoriesAS_0_dataarray_data_V_d0        => AS_D5PHIDn1_din
  );

  LATCH_TP_L1L2A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2A_bx,
      start => TP_L1L2A_start
  );

  TP_L1L2A : entity work.TP_L1L2A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => TP_done,
      bx_V          => TP_L1L2A_bx,
      bx_o_V        => TP_bx_out,
      bx_o_V_ap_vld => TP_bx_out_vld,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIA_BF_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIA_BF_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIA_BF_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIA_BF_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIA_BF_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIA_B_L1A_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIA_B_L1A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIA_B_L1A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIAn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIAn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIAn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIAn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIAn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIAn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIAn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIAn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIAn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIAn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIAn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIAn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIAn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIAn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIAn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIAn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIAn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIAn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIAn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIAn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIAn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIAn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIAn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIAn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2A_din
  );

  LATCH_TP_L1L2B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2B_bx,
      start => TP_L1L2B_start
  );

  TP_L1L2B : entity work.TP_L1L2B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIA_BE_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIA_BE_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIA_BE_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIA_BE_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIA_BE_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIB_BD_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIB_BD_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIB_BD_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIB_BD_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIB_BD_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIA_B_L1B_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIA_B_L1B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIA_B_L1B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIAn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIAn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIAn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIAn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIAn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIAn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIAn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIAn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIAn2_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIAn2_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIAn2_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIAn2_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIAn2_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIAn2_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIAn2_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIAn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIAn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIAn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIAn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIAn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIAn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIAn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIAn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIAn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2B_din
  );

  LATCH_TP_L1L2C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2C_bx,
      start => TP_L1L2C_start
  );

  TP_L1L2C : entity work.TP_L1L2C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIB_BC_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIB_BC_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIB_BC_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIB_BC_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIB_BC_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIC_BB_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIC_BB_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIC_BB_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIC_BB_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIC_BB_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIA_B_L1C_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIA_B_L1C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIA_B_L1C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIAn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIAn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIAn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIAn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIAn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIAn3_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIAn3_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIAn3_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIAn3_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIAn3_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIAn3_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIAn3_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIAn3_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIAn3_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIAn3_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIAn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIAn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIAn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIAn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIAn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIAn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIAn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIAn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIAn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2C_din
  );

  LATCH_TP_L1L2D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2D_bx,
      start => TP_L1L2D_start
  );

  TP_L1L2D : entity work.TP_L1L2D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIB_BA_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIB_BA_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIB_BA_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIB_BA_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIB_BA_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIC_BF_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIC_BF_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIC_BF_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIC_BF_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIC_BF_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIB_B_L1D_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIB_B_L1D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIB_B_L1D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIBn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIBn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIBn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIBn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIBn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIBn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIBn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIBn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIBn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIBn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIBn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIBn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIBn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIBn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIBn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIBn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIBn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIBn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIBn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIBn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIBn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIBn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIBn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIBn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2D_din
  );

  LATCH_TP_L1L2E: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2E_bx,
      start => TP_L1L2E_start
  );

  TP_L1L2E : entity work.TP_L1L2E
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2E_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2E_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIC_BE_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIC_BE_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIC_BE_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIC_BE_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIC_BE_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHID_BD_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHID_BD_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHID_BD_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHID_BD_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHID_BD_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIB_B_L1E_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIB_B_L1E_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIB_B_L1E_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIBn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIBn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIBn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIBn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIBn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIBn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIBn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIBn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIBn2_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIBn2_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIBn2_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIBn2_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIBn2_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIBn2_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIBn2_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIBn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIBn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIBn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIBn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIBn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIBn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIBn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIBn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIBn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2E_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2E_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2E_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2E_din
  );

  LATCH_TP_L1L2F: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2F_bx,
      start => TP_L1L2F_start
  );

  TP_L1L2F : entity work.TP_L1L2F
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2F_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2F_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHID_BC_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHID_BC_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHID_BC_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHID_BC_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHID_BC_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIE_BB_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIE_BB_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIE_BB_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIE_BB_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIE_BB_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIB_B_L1F_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIB_B_L1F_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIB_B_L1F_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIBn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIBn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIBn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIBn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIBn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIBn3_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIBn3_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIBn3_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIBn3_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIBn3_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIBn3_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIBn3_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIBn3_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIBn3_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIBn3_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIBn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIBn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIBn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIBn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIBn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIBn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIBn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIBn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIBn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2F_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2F_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2F_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2F_din
  );

  LATCH_TP_L1L2G: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2G_bx,
      start => TP_L1L2G_start
  );

  TP_L1L2G : entity work.TP_L1L2G
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2G_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2G_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHID_BA_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHID_BA_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHID_BA_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHID_BA_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHID_BA_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIE_BF_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIE_BF_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIE_BF_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIE_BF_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIE_BF_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIC_B_L1G_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIC_B_L1G_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIC_B_L1G_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHICn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHICn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHICn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHICn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHICn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHICn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHICn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHICn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHICn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHICn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHICn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHICn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHICn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHICn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHICn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHICn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHICn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHICn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHICn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHICn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHICn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHICn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHICn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHICn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2G_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2G_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2G_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2G_din
  );

  LATCH_TP_L1L2H: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2H_bx,
      start => TP_L1L2H_start
  );

  TP_L1L2H : entity work.TP_L1L2H
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2H_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2H_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIE_BE_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIE_BE_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIE_BE_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIE_BE_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIE_BE_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIF_BD_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIF_BD_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIF_BD_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIF_BD_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIF_BD_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIC_B_L1H_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIC_B_L1H_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIC_B_L1H_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHICn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHICn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHICn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHICn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHICn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHICn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHICn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHICn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHICn2_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHICn2_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHICn2_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHICn2_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHICn2_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHICn2_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHICn2_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHICn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHICn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHICn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHICn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHICn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHICn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHICn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHICn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHICn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2H_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2H_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2H_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2H_din
  );

  LATCH_TP_L1L2I: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2I_bx,
      start => TP_L1L2I_start
  );

  TP_L1L2I : entity work.TP_L1L2I
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2I_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2I_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIF_BC_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIF_BC_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIF_BC_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIF_BC_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIF_BC_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIG_BB_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIG_BB_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIG_BB_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIG_BB_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIG_BB_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHIC_B_L1I_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHIC_B_L1I_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHIC_B_L1I_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHICn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHICn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHICn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHICn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHICn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHICn3_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHICn3_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHICn3_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHICn3_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHICn3_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHICn3_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHICn3_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHICn3_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHICn3_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHICn3_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHICn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHICn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHICn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHICn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHICn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHICn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHICn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHICn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHICn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2I_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2I_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2I_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2I_din
  );

  LATCH_TP_L1L2J: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2J_bx,
      start => TP_L1L2J_start
  );

  TP_L1L2J : entity work.TP_L1L2J
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2J_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2J_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIF_BA_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIF_BA_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIF_BA_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIF_BA_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIF_BA_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIG_BF_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIG_BF_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIG_BF_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIG_BF_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIG_BF_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHID_B_L1J_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHID_B_L1J_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHID_B_L1J_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIDn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIDn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIDn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIDn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIDn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIDn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIDn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIDn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIDn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIDn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIDn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIDn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIDn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIDn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIDn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIDn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIDn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIDn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIDn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIDn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIDn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIDn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIDn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIDn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2J_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2J_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2J_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2J_din
  );

  LATCH_TP_L1L2K: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2K_bx,
      start => TP_L1L2K_start
  );

  TP_L1L2K : entity work.TP_L1L2K
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2K_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2K_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIG_BE_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIG_BE_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIG_BE_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIG_BE_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIG_BE_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIH_BD_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIH_BD_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIH_BD_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIH_BD_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIH_BD_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHID_B_L1K_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHID_B_L1K_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHID_B_L1K_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIDn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIDn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIDn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIDn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIDn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIDn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIDn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIDn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIDn2_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIDn2_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIDn2_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIDn2_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIDn2_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIDn2_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIDn2_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIDn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIDn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIDn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIDn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIDn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIDn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIDn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIDn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIDn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2K_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2K_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2K_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2K_din
  );

  LATCH_TP_L1L2L: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1L2L_bx,
      start => TP_L1L2L_start
  );

  TP_L1L2L : entity work.TP_L1L2L
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1L2L_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1L2L_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIH_BC_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIH_BC_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIH_BC_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIH_BC_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIH_BC_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L2PHID_B_L1L_enb,
      outerStubs_dataarray_data_V_address0  => AS_L2PHID_B_L1L_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L2PHID_B_L1L_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L2PHIDn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L2PHIDn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L2PHIDn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L2PHIDn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L2PHIDn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L2PHIDn3_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L2PHIDn3_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L2PHIDn3_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L2PHIDn3_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L2PHIDn3_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L2PHIDn3_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L2PHIDn3_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L2PHIDn3_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L2PHIDn3_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L2PHIDn3_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L2PHIDn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L2PHIDn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L2PHIDn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L2PHIDn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L2PHIDn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L2PHIDn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L2PHIDn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L2PHIDn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L2PHIDn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1L2L_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1L2L_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1L2L_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1L2L_din
  );

  LATCH_TP_L2L3A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2L3A_bx,
      start => TP_L2L3A_start
  );

  TP_L2L3A : entity work.TP_L2L3A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2L3A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2L3A_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHIA_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHIA_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHIA_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHIA_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHIA_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L3PHIA_B_L2A_enb,
      outerStubs_dataarray_data_V_address0  => AS_L3PHIA_B_L2A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L3PHIA_B_L2A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L3PHIIn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L3PHIIn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L3PHIIn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L3PHIIn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L3PHIIn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L3PHIIn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_L3PHIIn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L3PHIIn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L3PHIIn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L3PHIIn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L3PHIIn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L3PHIIn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L3PHIIn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L3PHIIn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L3PHIIn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2L3A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2L3A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2L3A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2L3A_din
  );

  LATCH_TP_L2L3B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2L3B_bx,
      start => TP_L2L3B_start
  );

  TP_L2L3B : entity work.TP_L2L3B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2L3B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2L3B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHIB_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHIB_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHIB_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHIB_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHIB_BM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L2PHIC_BL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L2PHIC_BL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L2PHIC_BL_V_dout,
      innerStubs_1_nentries_0_V               => AS_L2PHIC_BL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L2PHIC_BL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L3PHIB_B_L2B_enb,
      outerStubs_dataarray_data_V_address0  => AS_L3PHIB_B_L2B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L3PHIB_B_L2B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L3PHIJn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L3PHIJn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L3PHIJn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L3PHIJn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L3PHIJn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L3PHIJn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_L3PHIJn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L3PHIJn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L3PHIJn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L3PHIJn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L3PHIJn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L3PHIJn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L3PHIJn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L3PHIJn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L3PHIJn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2L3B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2L3B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2L3B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2L3B_din
  );

  LATCH_TP_L2L3C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2L3C_bx,
      start => TP_L2L3C_start
  );

  TP_L2L3C : entity work.TP_L2L3C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2L3C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2L3C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHIB_BR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHIB_BR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHIB_BR_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHIB_BR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHIB_BR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L2PHIC_BM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L2PHIC_BM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L2PHIC_BM_V_dout,
      innerStubs_1_nentries_0_V               => AS_L2PHIC_BM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L2PHIC_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L3PHIC_B_L2C_enb,
      outerStubs_dataarray_data_V_address0  => AS_L3PHIC_B_L2C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L3PHIC_B_L2C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L3PHIKn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L3PHIKn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L3PHIKn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L3PHIKn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L3PHIKn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L3PHIKn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_L3PHIKn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L3PHIKn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L3PHIKn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L3PHIKn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L3PHIKn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L3PHIKn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L3PHIKn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L3PHIKn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L3PHIKn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2L3C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2L3C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2L3C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2L3C_din
  );

  LATCH_TP_L2L3D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2L3D_bx,
      start => TP_L2L3D_start
  );

  TP_L2L3D : entity work.TP_L2L3D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2L3D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2L3D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHID_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHID_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHID_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHID_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHID_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L3PHID_B_L2D_enb,
      outerStubs_dataarray_data_V_address0  => AS_L3PHID_B_L2D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L3PHID_B_L2D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L3PHILn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L3PHILn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L3PHILn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L3PHILn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L3PHILn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L3PHILn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_L3PHILn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L3PHILn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L3PHILn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L3PHILn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L3PHILn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L3PHILn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L3PHILn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L3PHILn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L3PHILn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2L3D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2L3D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2L3D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2L3D_din
  );

  LATCH_TP_L3L4A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L3L4A_bx,
      start => TP_L3L4A_start
  );

  TP_L3L4A : entity work.TP_L3L4A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L3L4A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L3L4A_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L3PHIA_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L3PHIA_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L3PHIA_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L3PHIA_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L3PHIA_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L4PHIA_B_L3A_enb,
      outerStubs_dataarray_data_V_address0  => AS_L4PHIA_B_L3A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L4PHIA_B_L3A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L4PHIAn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L4PHIAn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L4PHIAn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L4PHIAn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L4PHIAn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L4PHIAn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L4PHIAn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L4PHIAn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L4PHIAn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L4PHIAn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L4PHIAn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L4PHIAn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L4PHIAn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L4PHIAn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L4PHIAn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L4PHIAn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L4PHIAn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L4PHIAn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L4PHIAn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L4PHIAn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L4PHIAn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L4PHIAn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L4PHIAn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L4PHIAn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L3L4A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L3L4A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L3L4A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L3L4A_din
  );

  LATCH_TP_L3L4B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L3L4B_bx,
      start => TP_L3L4B_start
  );

  TP_L3L4B : entity work.TP_L3L4B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L3L4B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L3L4B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L3PHIB_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L3PHIB_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L3PHIB_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L3PHIB_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L3PHIB_BM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L3PHIC_BL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L3PHIC_BL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L3PHIC_BL_V_dout,
      innerStubs_1_nentries_0_V               => AS_L3PHIC_BL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L3PHIC_BL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L4PHIB_B_L3B_enb,
      outerStubs_dataarray_data_V_address0  => AS_L4PHIB_B_L3B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L4PHIB_B_L3B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L4PHIBn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L4PHIBn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L4PHIBn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L4PHIBn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L4PHIBn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L4PHIBn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L4PHIBn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L4PHIBn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L4PHIBn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L4PHIBn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L4PHIBn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L4PHIBn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L4PHIBn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L4PHIBn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L4PHIBn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L4PHIBn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L4PHIBn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L4PHIBn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L4PHIBn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L4PHIBn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L4PHIBn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L4PHIBn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L4PHIBn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L4PHIBn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L3L4B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L3L4B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L3L4B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L3L4B_din
  );

  LATCH_TP_L3L4C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L3L4C_bx,
      start => TP_L3L4C_start
  );

  TP_L3L4C : entity work.TP_L3L4C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L3L4C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L3L4C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L3PHIB_BR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L3PHIB_BR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L3PHIB_BR_V_dout,
      innerStubs_0_nentries_0_V               => AS_L3PHIB_BR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L3PHIB_BR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L3PHIC_BM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L3PHIC_BM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L3PHIC_BM_V_dout,
      innerStubs_1_nentries_0_V               => AS_L3PHIC_BM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L3PHIC_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L4PHIC_B_L3C_enb,
      outerStubs_dataarray_data_V_address0  => AS_L4PHIC_B_L3C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L4PHIC_B_L3C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L4PHICn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L4PHICn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L4PHICn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L4PHICn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L4PHICn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L4PHICn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L4PHICn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L4PHICn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L4PHICn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L4PHICn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L4PHICn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L4PHICn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L4PHICn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L4PHICn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L4PHICn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L4PHICn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L4PHICn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L4PHICn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L4PHICn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L4PHICn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L4PHICn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L4PHICn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L4PHICn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L4PHICn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L3L4C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L3L4C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L3L4C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L3L4C_din
  );

  LATCH_TP_L3L4D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L3L4D_bx,
      start => TP_L3L4D_start
  );

  TP_L3L4D : entity work.TP_L3L4D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L3L4D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L3L4D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L3PHID_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L3PHID_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L3PHID_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L3PHID_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L3PHID_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L4PHID_B_L3D_enb,
      outerStubs_dataarray_data_V_address0  => AS_L4PHID_B_L3D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L4PHID_B_L3D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L4PHIDn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L4PHIDn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L4PHIDn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L4PHIDn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L4PHIDn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L4PHIDn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L4PHIDn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L4PHIDn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L4PHIDn1_AV_dout(2),
      outerVMStubs_dataarray_3_data_V_ce0       => VMSTE_L4PHIDn1_A_enb(3),
      outerVMStubs_dataarray_3_data_V_address0  => VMSTE_L4PHIDn1_AV_readaddr(3),
      outerVMStubs_dataarray_3_data_V_q0        => VMSTE_L4PHIDn1_AV_dout(3),
      outerVMStubs_dataarray_4_data_V_ce0       => VMSTE_L4PHIDn1_A_enb(4),
      outerVMStubs_dataarray_4_data_V_address0  => VMSTE_L4PHIDn1_AV_readaddr(4),
      outerVMStubs_dataarray_4_data_V_q0        => VMSTE_L4PHIDn1_AV_dout(4),
      outerVMStubs_nentries_V_ce0 => VMSTE_L4PHIDn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L4PHIDn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L4PHIDn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L4PHIDn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L4PHIDn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L4PHIDn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L4PHIDn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L4PHIDn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L4PHIDn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L3L4D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L3L4D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L3L4D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L3L4D_din
  );

  LATCH_TP_L5L6A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L5L6A_bx,
      start => TP_L5L6A_start
  );

  TP_L5L6A : entity work.TP_L5L6A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L5L6A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L5L6A_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L5PHIA_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L5PHIA_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L5PHIA_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L5PHIA_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L5PHIA_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L6PHIA_B_L5A_enb,
      outerStubs_dataarray_data_V_address0  => AS_L6PHIA_B_L5A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L6PHIA_B_L5A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L6PHIAn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L6PHIAn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L6PHIAn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L6PHIAn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L6PHIAn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L6PHIAn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L6PHIAn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L6PHIAn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L6PHIAn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_L6PHIAn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L6PHIAn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L6PHIAn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L6PHIAn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L6PHIAn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L6PHIAn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L6PHIAn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L6PHIAn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L6PHIAn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L5L6A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L5L6A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L5L6A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L5L6A_din
  );

  LATCH_TP_L5L6B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L5L6B_bx,
      start => TP_L5L6B_start
  );

  TP_L5L6B : entity work.TP_L5L6B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L5L6B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L5L6B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L5PHIB_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L5PHIB_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L5PHIB_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L5PHIB_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L5PHIB_BM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L5PHIC_BL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L5PHIC_BL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L5PHIC_BL_V_dout,
      innerStubs_1_nentries_0_V               => AS_L5PHIC_BL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L5PHIC_BL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L6PHIB_B_L5B_enb,
      outerStubs_dataarray_data_V_address0  => AS_L6PHIB_B_L5B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L6PHIB_B_L5B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L6PHIBn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L6PHIBn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L6PHIBn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L6PHIBn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L6PHIBn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L6PHIBn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L6PHIBn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L6PHIBn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L6PHIBn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_L6PHIBn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L6PHIBn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L6PHIBn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L6PHIBn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L6PHIBn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L6PHIBn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L6PHIBn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L6PHIBn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L6PHIBn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L5L6B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L5L6B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L5L6B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L5L6B_din
  );

  LATCH_TP_L5L6C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L5L6C_bx,
      start => TP_L5L6C_start
  );

  TP_L5L6C : entity work.TP_L5L6C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L5L6C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L5L6C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L5PHIB_BR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L5PHIB_BR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L5PHIB_BR_V_dout,
      innerStubs_0_nentries_0_V               => AS_L5PHIB_BR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L5PHIB_BR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L5PHIC_BM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L5PHIC_BM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L5PHIC_BM_V_dout,
      innerStubs_1_nentries_0_V               => AS_L5PHIC_BM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L5PHIC_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L6PHIC_B_L5C_enb,
      outerStubs_dataarray_data_V_address0  => AS_L6PHIC_B_L5C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L6PHIC_B_L5C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L6PHICn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L6PHICn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L6PHICn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L6PHICn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L6PHICn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L6PHICn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L6PHICn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L6PHICn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L6PHICn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_L6PHICn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L6PHICn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L6PHICn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L6PHICn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L6PHICn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L6PHICn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L6PHICn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L6PHICn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L6PHICn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L5L6C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L5L6C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L5L6C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L5L6C_din
  );

  LATCH_TP_L5L6D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L5L6D_bx,
      start => TP_L5L6D_start
  );

  TP_L5L6D : entity work.TP_L5L6D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L5L6D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L5L6D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L5PHID_BM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L5PHID_BM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L5PHID_BM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L5PHID_BM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L5PHID_BM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_L6PHID_B_L5D_enb,
      outerStubs_dataarray_data_V_address0  => AS_L6PHID_B_L5D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_L6PHID_B_L5D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_L6PHIDn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_L6PHIDn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_L6PHIDn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_L6PHIDn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_L6PHIDn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_L6PHIDn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_L6PHIDn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_L6PHIDn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_L6PHIDn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_L6PHIDn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_L6PHIDn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_L6PHIDn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_L6PHIDn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_L6PHIDn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_L6PHIDn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_L6PHIDn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_L6PHIDn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_L6PHIDn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L5L6D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L5L6D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L5L6D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L5L6D_din
  );

  LATCH_TP_D1D2A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D1D2A_bx,
      start => TP_D1D2A_start
  );

  TP_D1D2A : entity work.TP_D1D2A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D1D2A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D1D2A_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D1PHIA_DM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D1PHIA_DM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D1PHIA_DM_V_dout,
      innerStubs_0_nentries_0_V               => AS_D1PHIA_DM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D1PHIA_DM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D2PHIA_D_D1A_enb,
      outerStubs_dataarray_data_V_address0  => AS_D2PHIA_D_D1A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D2PHIA_D_D1A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D2PHIAn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D2PHIAn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D2PHIAn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D2PHIAn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D2PHIAn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D2PHIAn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D2PHIAn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D2PHIAn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D2PHIAn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D2PHIAn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D2PHIAn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D2PHIAn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D2PHIAn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D2PHIAn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D2PHIAn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D2PHIAn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D2PHIAn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D2PHIAn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D1D2A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D1D2A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D1D2A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D1D2A_din
  );

  LATCH_TP_D1D2B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D1D2B_bx,
      start => TP_D1D2B_start
  );

  TP_D1D2B : entity work.TP_D1D2B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D1D2B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D1D2B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D1PHIB_DM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D1PHIB_DM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D1PHIB_DM_V_dout,
      innerStubs_0_nentries_0_V               => AS_D1PHIB_DM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D1PHIB_DM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_D1PHIC_DL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_D1PHIC_DL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_D1PHIC_DL_V_dout,
      innerStubs_1_nentries_0_V               => AS_D1PHIC_DL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_D1PHIC_DL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D2PHIB_D_D1B_enb,
      outerStubs_dataarray_data_V_address0  => AS_D2PHIB_D_D1B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D2PHIB_D_D1B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D2PHIBn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D2PHIBn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D2PHIBn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D2PHIBn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D2PHIBn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D2PHIBn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D2PHIBn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D2PHIBn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D2PHIBn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D2PHIBn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D2PHIBn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D2PHIBn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D2PHIBn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D2PHIBn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D2PHIBn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D2PHIBn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D2PHIBn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D2PHIBn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D1D2B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D1D2B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D1D2B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D1D2B_din
  );

  LATCH_TP_D1D2C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D1D2C_bx,
      start => TP_D1D2C_start
  );

  TP_D1D2C : entity work.TP_D1D2C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D1D2C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D1D2C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D1PHIB_DR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D1PHIB_DR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D1PHIB_DR_V_dout,
      innerStubs_0_nentries_0_V               => AS_D1PHIB_DR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D1PHIB_DR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_D1PHIC_DM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_D1PHIC_DM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_D1PHIC_DM_V_dout,
      innerStubs_1_nentries_0_V               => AS_D1PHIC_DM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_D1PHIC_DM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D2PHIC_D_D1C_enb,
      outerStubs_dataarray_data_V_address0  => AS_D2PHIC_D_D1C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D2PHIC_D_D1C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D2PHICn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D2PHICn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D2PHICn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D2PHICn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D2PHICn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D2PHICn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D2PHICn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D2PHICn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D2PHICn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D2PHICn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D2PHICn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D2PHICn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D2PHICn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D2PHICn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D2PHICn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D2PHICn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D2PHICn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D2PHICn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D1D2C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D1D2C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D1D2C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D1D2C_din
  );

  LATCH_TP_D1D2D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D1D2D_bx,
      start => TP_D1D2D_start
  );

  TP_D1D2D : entity work.TP_D1D2D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D1D2D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D1D2D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D1PHID_DM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D1PHID_DM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D1PHID_DM_V_dout,
      innerStubs_0_nentries_0_V               => AS_D1PHID_DM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D1PHID_DM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D2PHID_D_D1D_enb,
      outerStubs_dataarray_data_V_address0  => AS_D2PHID_D_D1D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D2PHID_D_D1D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D2PHIDn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D2PHIDn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D2PHIDn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D2PHIDn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D2PHIDn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D2PHIDn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D2PHIDn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D2PHIDn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D2PHIDn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D2PHIDn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D2PHIDn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D2PHIDn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D2PHIDn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D2PHIDn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D2PHIDn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D2PHIDn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D2PHIDn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D2PHIDn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D1D2D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D1D2D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D1D2D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D1D2D_din
  );

  LATCH_TP_D3D4A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D3D4A_bx,
      start => TP_D3D4A_start
  );

  TP_D3D4A : entity work.TP_D3D4A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D3D4A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D3D4A_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D3PHIA_DM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D3PHIA_DM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D3PHIA_DM_V_dout,
      innerStubs_0_nentries_0_V               => AS_D3PHIA_DM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D3PHIA_DM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D4PHIA_D_D3A_enb,
      outerStubs_dataarray_data_V_address0  => AS_D4PHIA_D_D3A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D4PHIA_D_D3A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D4PHIAn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D4PHIAn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D4PHIAn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D4PHIAn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D4PHIAn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D4PHIAn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D4PHIAn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D4PHIAn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D4PHIAn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D4PHIAn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D4PHIAn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D4PHIAn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D4PHIAn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D4PHIAn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D4PHIAn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D3D4A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D3D4A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D3D4A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D3D4A_din
  );

  LATCH_TP_D3D4B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D3D4B_bx,
      start => TP_D3D4B_start
  );

  TP_D3D4B : entity work.TP_D3D4B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D3D4B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D3D4B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D3PHIB_DM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D3PHIB_DM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D3PHIB_DM_V_dout,
      innerStubs_0_nentries_0_V               => AS_D3PHIB_DM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D3PHIB_DM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_D3PHIC_DL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_D3PHIC_DL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_D3PHIC_DL_V_dout,
      innerStubs_1_nentries_0_V               => AS_D3PHIC_DL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_D3PHIC_DL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D4PHIB_D_D3B_enb,
      outerStubs_dataarray_data_V_address0  => AS_D4PHIB_D_D3B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D4PHIB_D_D3B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D4PHIBn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D4PHIBn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D4PHIBn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D4PHIBn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D4PHIBn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D4PHIBn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D4PHIBn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D4PHIBn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D4PHIBn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D4PHIBn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D4PHIBn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D4PHIBn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D4PHIBn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D4PHIBn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D4PHIBn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D3D4B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D3D4B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D3D4B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D3D4B_din
  );

  LATCH_TP_D3D4C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D3D4C_bx,
      start => TP_D3D4C_start
  );

  TP_D3D4C : entity work.TP_D3D4C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D3D4C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D3D4C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D3PHIB_DR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D3PHIB_DR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D3PHIB_DR_V_dout,
      innerStubs_0_nentries_0_V               => AS_D3PHIB_DR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D3PHIB_DR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_D3PHIC_DM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_D3PHIC_DM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_D3PHIC_DM_V_dout,
      innerStubs_1_nentries_0_V               => AS_D3PHIC_DM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_D3PHIC_DM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D4PHIC_D_D3C_enb,
      outerStubs_dataarray_data_V_address0  => AS_D4PHIC_D_D3C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D4PHIC_D_D3C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D4PHICn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D4PHICn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D4PHICn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D4PHICn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D4PHICn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D4PHICn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D4PHICn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D4PHICn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D4PHICn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D4PHICn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D4PHICn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D4PHICn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D4PHICn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D4PHICn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D4PHICn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D3D4C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D3D4C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D3D4C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D3D4C_din
  );

  LATCH_TP_D3D4D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_D3D4D_bx,
      start => TP_D3D4D_start
  );

  TP_D3D4D : entity work.TP_D3D4D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_D3D4D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_D3D4D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_D3PHID_DM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_D3PHID_DM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_D3PHID_DM_V_dout,
      innerStubs_0_nentries_0_V               => AS_D3PHID_DM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_D3PHID_DM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D4PHID_D_D3D_enb,
      outerStubs_dataarray_data_V_address0  => AS_D4PHID_D_D3D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D4PHID_D_D3D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D4PHIDn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D4PHIDn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D4PHIDn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D4PHIDn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D4PHIDn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D4PHIDn1_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D4PHIDn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D4PHIDn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D4PHIDn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D4PHIDn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D4PHIDn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D4PHIDn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D4PHIDn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D4PHIDn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D4PHIDn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_D3D4D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_D3D4D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_D3D4D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_D3D4D_din
  );

  LATCH_TP_L1D1A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1A_bx,
      start => TP_L1D1A_start
  );

  TP_L1D1A : entity work.TP_L1D1A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1A_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIA_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIA_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIA_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIA_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIA_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIA_O_L1A_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIA_O_L1A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIA_O_L1A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIXn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIXn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIXn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIXn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIXn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIXn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIXn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIXn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIXn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIXn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIXn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIXn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIXn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIXn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIXn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIXn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIXn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIXn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1A_din
  );

  LATCH_TP_L1D1B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1B_bx,
      start => TP_L1D1B_start
  );

  TP_L1D1B : entity work.TP_L1D1B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIB_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIB_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIB_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIB_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIB_OM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIC_OL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIC_OL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIC_OL_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIC_OL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIC_OL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIA_O_L1B_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIA_O_L1B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIA_O_L1B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIXn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIXn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIXn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIXn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIXn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIXn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIXn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIXn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIXn2_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIXn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIXn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIXn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIXn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIXn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIXn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIXn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIXn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIXn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1B_din
  );

  LATCH_TP_L1D1C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1C_bx,
      start => TP_L1D1C_start
  );

  TP_L1D1C : entity work.TP_L1D1C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIB_OR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIB_OR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIB_OR_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIB_OR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIB_OR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIC_OM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIC_OM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIC_OM_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIC_OM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIC_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIB_O_L1C_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIB_O_L1C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIB_O_L1C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIYn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIYn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIYn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIYn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIYn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIYn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIYn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIYn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIYn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIYn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIYn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIYn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIYn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIYn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIYn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIYn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIYn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIYn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1C_din
  );

  LATCH_TP_L1D1D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1D_bx,
      start => TP_L1D1D_start
  );

  TP_L1D1D : entity work.TP_L1D1D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHID_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHID_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHID_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHID_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHID_OM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIE_OL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIE_OL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIE_OL_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIE_OL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIE_OL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIB_O_L1D_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIB_O_L1D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIB_O_L1D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIYn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIYn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIYn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIYn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIYn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIYn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIYn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIYn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIYn2_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIYn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIYn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIYn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIYn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIYn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIYn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIYn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIYn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIYn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1D_din
  );

  LATCH_TP_L1D1E: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1E_bx,
      start => TP_L1D1E_start
  );

  TP_L1D1E : entity work.TP_L1D1E
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1E_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1E_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHID_OR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHID_OR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHID_OR_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHID_OR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHID_OR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIE_OM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIE_OM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIE_OM_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIE_OM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIE_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIC_O_L1E_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIC_O_L1E_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIC_O_L1E_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIZn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIZn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIZn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIZn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIZn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIZn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIZn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIZn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIZn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIZn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIZn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIZn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIZn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIZn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIZn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIZn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIZn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIZn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1E_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1E_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1E_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1E_din
  );

  LATCH_TP_L1D1F: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1F_bx,
      start => TP_L1D1F_start
  );

  TP_L1D1F : entity work.TP_L1D1F
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1F_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1F_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIF_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIF_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIF_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIF_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIF_OM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIG_OL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIG_OL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIG_OL_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIG_OL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIG_OL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIC_O_L1F_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIC_O_L1F_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIC_O_L1F_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIZn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIZn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIZn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIZn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIZn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIZn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIZn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIZn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIZn2_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIZn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIZn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIZn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIZn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIZn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIZn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIZn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIZn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIZn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1F_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1F_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1F_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1F_din
  );

  LATCH_TP_L1D1G: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1G_bx,
      start => TP_L1D1G_start
  );

  TP_L1D1G : entity work.TP_L1D1G
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1G_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1G_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIF_OR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIF_OR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIF_OR_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIF_OR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIF_OR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L1PHIG_OM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L1PHIG_OM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L1PHIG_OM_V_dout,
      innerStubs_1_nentries_0_V               => AS_L1PHIG_OM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L1PHIG_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHID_O_L1G_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHID_O_L1G_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHID_O_L1G_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIWn1_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIWn1_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIWn1_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIWn1_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIWn1_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIWn1_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIWn1_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIWn1_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIWn1_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIWn1_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIWn1_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIWn1_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIWn1_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIWn1_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIWn1_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIWn1_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIWn1_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIWn1_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1G_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1G_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1G_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1G_din
  );

  LATCH_TP_L1D1H: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L1D1H_bx,
      start => TP_L1D1H_start
  );

  TP_L1D1H : entity work.TP_L1D1H
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L1D1H_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L1D1H_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L1PHIH_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L1PHIH_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L1PHIH_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L1PHIH_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L1PHIH_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHID_O_L1H_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHID_O_L1H_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHID_O_L1H_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIWn2_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIWn2_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIWn2_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIWn2_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIWn2_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIWn2_AV_dout(1),
      outerVMStubs_dataarray_2_data_V_ce0       => VMSTE_D1PHIWn2_A_enb(2),
      outerVMStubs_dataarray_2_data_V_address0  => VMSTE_D1PHIWn2_AV_readaddr(2),
      outerVMStubs_dataarray_2_data_V_q0        => VMSTE_D1PHIWn2_AV_dout(2),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIWn2_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIWn2_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIWn2_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIWn2_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIWn2_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIWn2_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIWn2_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIWn2_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIWn2_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L1D1H_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L1D1H_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L1D1H_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L1D1H_din
  );

  LATCH_TP_L2D1A: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2D1A_bx,
      start => TP_L2D1A_start
  );

  TP_L2D1A : entity work.TP_L2D1A
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2D1A_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2D1A_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHIA_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHIA_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHIA_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHIA_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHIA_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIA_O_L2A_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIA_O_L2A_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIA_O_L2A_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIXn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIXn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIXn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIXn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIXn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIXn3_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIXn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIXn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIXn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIXn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIXn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIXn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIXn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIXn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIXn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2D1A_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2D1A_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2D1A_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2D1A_din
  );

  LATCH_TP_L2D1B: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2D1B_bx,
      start => TP_L2D1B_start
  );

  TP_L2D1B : entity work.TP_L2D1B
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2D1B_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2D1B_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHIB_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHIB_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHIB_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHIB_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHIB_OM_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L2PHIC_OL_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L2PHIC_OL_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L2PHIC_OL_V_dout,
      innerStubs_1_nentries_0_V               => AS_L2PHIC_OL_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L2PHIC_OL_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIB_O_L2B_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIB_O_L2B_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIB_O_L2B_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIYn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIYn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIYn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIYn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIYn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIYn3_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIYn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIYn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIYn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIYn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIYn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIYn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIYn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIYn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIYn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2D1B_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2D1B_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2D1B_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2D1B_din
  );

  LATCH_TP_L2D1C: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2D1C_bx,
      start => TP_L2D1C_start
  );

  TP_L2D1C : entity work.TP_L2D1C
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2D1C_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2D1C_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHIB_OR_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHIB_OR_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHIB_OR_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHIB_OR_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHIB_OR_AV_dout_nent(1),
      innerStubs_1_dataarray_data_V_ce0       => AS_L2PHIC_OM_enb,
      innerStubs_1_dataarray_data_V_address0  => AS_L2PHIC_OM_V_readaddr,
      innerStubs_1_dataarray_data_V_q0        => AS_L2PHIC_OM_V_dout,
      innerStubs_1_nentries_0_V               => AS_L2PHIC_OM_AV_dout_nent(0),
      innerStubs_1_nentries_1_V               => AS_L2PHIC_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHIC_O_L2C_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHIC_O_L2C_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHIC_O_L2C_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIZn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIZn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIZn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIZn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIZn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIZn3_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIZn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIZn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIZn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIZn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIZn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIZn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIZn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIZn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIZn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2D1C_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2D1C_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2D1C_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2D1C_din
  );

  LATCH_TP_L2D1D: entity work.tf_pipeline_slr_xing
    port map (
      clk   => clk,
      done  => VMR_done,
      bx_out => VMR_bx_out,
      bx => TP_L2D1D_bx,
      start => TP_L2D1D_start
  );

  TP_L2D1D : entity work.TP_L2D1D
    port map (
      ap_clk   => clk,
      ap_rst   => reset,
      ap_start => TP_L2D1D_start,
      ap_idle  => open,
      ap_ready => open,
      ap_done  => open,
      bx_V          => TP_L2D1D_bx,
      innerStubs_0_dataarray_data_V_ce0       => AS_L2PHID_OM_enb,
      innerStubs_0_dataarray_data_V_address0  => AS_L2PHID_OM_V_readaddr,
      innerStubs_0_dataarray_data_V_q0        => AS_L2PHID_OM_V_dout,
      innerStubs_0_nentries_0_V               => AS_L2PHID_OM_AV_dout_nent(0),
      innerStubs_0_nentries_1_V               => AS_L2PHID_OM_AV_dout_nent(1),
      outerStubs_dataarray_data_V_ce0       => AS_D1PHID_O_L2D_enb,
      outerStubs_dataarray_data_V_address0  => AS_D1PHID_O_L2D_V_readaddr,
      outerStubs_dataarray_data_V_q0        => AS_D1PHID_O_L2D_V_dout,
      outerVMStubs_dataarray_0_data_V_ce0       => VMSTE_D1PHIWn3_A_enb(0),
      outerVMStubs_dataarray_0_data_V_address0  => VMSTE_D1PHIWn3_AV_readaddr(0),
      outerVMStubs_dataarray_0_data_V_q0        => VMSTE_D1PHIWn3_AV_dout(0),
      outerVMStubs_dataarray_1_data_V_ce0       => VMSTE_D1PHIWn3_A_enb(1),
      outerVMStubs_dataarray_1_data_V_address0  => VMSTE_D1PHIWn3_AV_readaddr(1),
      outerVMStubs_dataarray_1_data_V_q0        => VMSTE_D1PHIWn3_AV_dout(1),
      outerVMStubs_nentries_V_ce0 => VMSTE_D1PHIWn3_enb_nent,
      outerVMStubs_nentries_V_address0 => VMSTE_D1PHIWn3_V_addr_nent,
      outerVMStubs_nentries_V_q0 => VMSTE_D1PHIWn3_AV_dout_nent,
      outerVMStubs_binmaskA_V_address0 => VMSTE_D1PHIWn3_V_addr_binmaskA,
      outerVMStubs_binmaskA_V_ce0 => VMSTE_D1PHIWn3_enb_binmaskA,
      outerVMStubs_binmaskA_V_q0 => VMSTE_D1PHIWn3_V_binmaskA,
      outerVMStubs_binmaskB_V_address0 => VMSTE_D1PHIWn3_V_addr_binmaskB,
      outerVMStubs_binmaskB_V_ce0 => VMSTE_D1PHIWn3_enb_binmaskB,
      outerVMStubs_binmaskB_V_q0 => VMSTE_D1PHIWn3_V_binmaskB,
      trackletParameters_dataarray_data_V_ce0       => open,
      trackletParameters_dataarray_data_V_we0       => TPAR_L2D1D_wea,
      trackletParameters_dataarray_data_V_address0(9 downto 0)  => TPAR_L2D1D_writeaddr,
      trackletParameters_dataarray_data_V_address0(11 downto 10)  => TPAR_L2D1D_dummy,
      trackletParameters_dataarray_data_V_d0        => TPAR_L2D1D_din
  );

end rtl;
